`ifdef ST_WIDTH_INF_16
$fwrite(tri_report_ieee754, "===============================%d Column Results    ======================================\n",col_index);
$fwrite(tri_report_ieee754, "Item0   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent0  , golden_yjp0  , dut_yjp0  );
$fwrite(tri_report_ieee754, "Item1   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent1  , golden_yjp1  , dut_yjp1  );
$fwrite(tri_report_ieee754, "Item2   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent2  , golden_yjp2  , dut_yjp2  );
$fwrite(tri_report_ieee754, "Item3   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent3  , golden_yjp3  , dut_yjp3  );
$fwrite(tri_report_ieee754, "Item4   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent4  , golden_yjp4  , dut_yjp4  );
$fwrite(tri_report_ieee754, "Item5   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent5  , golden_yjp5  , dut_yjp5  );
$fwrite(tri_report_ieee754, "Item6   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent6  , golden_yjp6  , dut_yjp6  );
$fwrite(tri_report_ieee754, "Item7   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent7  , golden_yjp7  , dut_yjp7  );
`endif // ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_256
$fwrite(tri_report_ieee754, "Item8   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent8  , golden_yjp8  , dut_yjp8  );
$fwrite(tri_report_ieee754, "Item9   error percent: %f%%, golden result: %h, dut result: %h\n", error_percent9  , golden_yjp9  , dut_yjp9  );
$fwrite(tri_report_ieee754, "Item10  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent10 , golden_yjp10 , dut_yjp10 );
$fwrite(tri_report_ieee754, "Item11  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent11 , golden_yjp11 , dut_yjp11 );
$fwrite(tri_report_ieee754, "Item12  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent12 , golden_yjp12 , dut_yjp12 );
$fwrite(tri_report_ieee754, "Item13  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent13 , golden_yjp13 , dut_yjp13 );
$fwrite(tri_report_ieee754, "Item14  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent14 , golden_yjp14 , dut_yjp14 );
$fwrite(tri_report_ieee754, "Item15  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent15 , golden_yjp15 , dut_yjp15 );
$fwrite(tri_report_ieee754, "Item16  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent16 , golden_yjp16 , dut_yjp16 );
$fwrite(tri_report_ieee754, "Item17  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent17 , golden_yjp17 , dut_yjp17 );
$fwrite(tri_report_ieee754, "Item18  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent18 , golden_yjp18 , dut_yjp18 );
$fwrite(tri_report_ieee754, "Item19  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent19 , golden_yjp19 , dut_yjp19 );
$fwrite(tri_report_ieee754, "Item20  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent20 , golden_yjp20 , dut_yjp20 );
$fwrite(tri_report_ieee754, "Item21  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent21 , golden_yjp21 , dut_yjp21 );
$fwrite(tri_report_ieee754, "Item22  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent22 , golden_yjp22 , dut_yjp22 );
$fwrite(tri_report_ieee754, "Item23  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent23 , golden_yjp23 , dut_yjp23 );
$fwrite(tri_report_ieee754, "Item24  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent24 , golden_yjp24 , dut_yjp24 );
$fwrite(tri_report_ieee754, "Item25  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent25 , golden_yjp25 , dut_yjp25 );
$fwrite(tri_report_ieee754, "Item26  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent26 , golden_yjp26 , dut_yjp26 );
$fwrite(tri_report_ieee754, "Item27  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent27 , golden_yjp27 , dut_yjp27 );
$fwrite(tri_report_ieee754, "Item28  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent28 , golden_yjp28 , dut_yjp28 );
$fwrite(tri_report_ieee754, "Item29  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent29 , golden_yjp29 , dut_yjp29 );
$fwrite(tri_report_ieee754, "Item30  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent30 , golden_yjp30 , dut_yjp30 );
$fwrite(tri_report_ieee754, "Item31  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent31 , golden_yjp31 , dut_yjp31 );
$fwrite(tri_report_ieee754, "Item32  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent32 , golden_yjp32 , dut_yjp32 );
$fwrite(tri_report_ieee754, "Item33  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent33 , golden_yjp33 , dut_yjp33 );
$fwrite(tri_report_ieee754, "Item34  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent34 , golden_yjp34 , dut_yjp34 );
$fwrite(tri_report_ieee754, "Item35  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent35 , golden_yjp35 , dut_yjp35 );
$fwrite(tri_report_ieee754, "Item36  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent36 , golden_yjp36 , dut_yjp36 );
$fwrite(tri_report_ieee754, "Item37  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent37 , golden_yjp37 , dut_yjp37 );
$fwrite(tri_report_ieee754, "Item38  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent38 , golden_yjp38 , dut_yjp38 );
$fwrite(tri_report_ieee754, "Item39  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent39 , golden_yjp39 , dut_yjp39 );
$fwrite(tri_report_ieee754, "Item40  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent40 , golden_yjp40 , dut_yjp40 );
$fwrite(tri_report_ieee754, "Item41  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent41 , golden_yjp41 , dut_yjp41 );
$fwrite(tri_report_ieee754, "Item42  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent42 , golden_yjp42 , dut_yjp42 );
$fwrite(tri_report_ieee754, "Item43  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent43 , golden_yjp43 , dut_yjp43 );
$fwrite(tri_report_ieee754, "Item44  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent44 , golden_yjp44 , dut_yjp44 );
$fwrite(tri_report_ieee754, "Item45  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent45 , golden_yjp45 , dut_yjp45 );
$fwrite(tri_report_ieee754, "Item46  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent46 , golden_yjp46 , dut_yjp46 );
$fwrite(tri_report_ieee754, "Item47  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent47 , golden_yjp47 , dut_yjp47 );
$fwrite(tri_report_ieee754, "Item48  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent48 , golden_yjp48 , dut_yjp48 );
$fwrite(tri_report_ieee754, "Item49  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent49 , golden_yjp49 , dut_yjp49 );
$fwrite(tri_report_ieee754, "Item50  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent50 , golden_yjp50 , dut_yjp50 );
$fwrite(tri_report_ieee754, "Item51  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent51 , golden_yjp51 , dut_yjp51 );
$fwrite(tri_report_ieee754, "Item52  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent52 , golden_yjp52 , dut_yjp52 );
$fwrite(tri_report_ieee754, "Item53  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent53 , golden_yjp53 , dut_yjp53 );
$fwrite(tri_report_ieee754, "Item54  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent54 , golden_yjp54 , dut_yjp54 );
$fwrite(tri_report_ieee754, "Item55  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent55 , golden_yjp55 , dut_yjp55 );
$fwrite(tri_report_ieee754, "Item56  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent56 , golden_yjp56 , dut_yjp56 );
$fwrite(tri_report_ieee754, "Item57  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent57 , golden_yjp57 , dut_yjp57 );
$fwrite(tri_report_ieee754, "Item58  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent58 , golden_yjp58 , dut_yjp58 );
$fwrite(tri_report_ieee754, "Item59  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent59 , golden_yjp59 , dut_yjp59 );
$fwrite(tri_report_ieee754, "Item60  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent60 , golden_yjp60 , dut_yjp60 );
$fwrite(tri_report_ieee754, "Item61  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent61 , golden_yjp61 , dut_yjp61 );
$fwrite(tri_report_ieee754, "Item62  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent62 , golden_yjp62 , dut_yjp62 );
$fwrite(tri_report_ieee754, "Item63  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent63 , golden_yjp63 , dut_yjp63 );
$fwrite(tri_report_ieee754, "Item64  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent64 , golden_yjp64 , dut_yjp64 );
$fwrite(tri_report_ieee754, "Item65  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent65 , golden_yjp65 , dut_yjp65 );
$fwrite(tri_report_ieee754, "Item66  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent66 , golden_yjp66 , dut_yjp66 );
$fwrite(tri_report_ieee754, "Item67  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent67 , golden_yjp67 , dut_yjp67 );
$fwrite(tri_report_ieee754, "Item68  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent68 , golden_yjp68 , dut_yjp68 );
$fwrite(tri_report_ieee754, "Item69  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent69 , golden_yjp69 , dut_yjp69 );
$fwrite(tri_report_ieee754, "Item70  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent70 , golden_yjp70 , dut_yjp70 );
$fwrite(tri_report_ieee754, "Item71  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent71 , golden_yjp71 , dut_yjp71 );
$fwrite(tri_report_ieee754, "Item72  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent72 , golden_yjp72 , dut_yjp72 );
$fwrite(tri_report_ieee754, "Item73  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent73 , golden_yjp73 , dut_yjp73 );
$fwrite(tri_report_ieee754, "Item74  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent74 , golden_yjp74 , dut_yjp74 );
$fwrite(tri_report_ieee754, "Item75  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent75 , golden_yjp75 , dut_yjp75 );
$fwrite(tri_report_ieee754, "Item76  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent76 , golden_yjp76 , dut_yjp76 );
$fwrite(tri_report_ieee754, "Item77  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent77 , golden_yjp77 , dut_yjp77 );
$fwrite(tri_report_ieee754, "Item78  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent78 , golden_yjp78 , dut_yjp78 );
$fwrite(tri_report_ieee754, "Item79  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent79 , golden_yjp79 , dut_yjp79 );
$fwrite(tri_report_ieee754, "Item80  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent80 , golden_yjp80 , dut_yjp80 );
$fwrite(tri_report_ieee754, "Item81  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent81 , golden_yjp81 , dut_yjp81 );
$fwrite(tri_report_ieee754, "Item82  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent82 , golden_yjp82 , dut_yjp82 );
$fwrite(tri_report_ieee754, "Item83  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent83 , golden_yjp83 , dut_yjp83 );
$fwrite(tri_report_ieee754, "Item84  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent84 , golden_yjp84 , dut_yjp84 );
$fwrite(tri_report_ieee754, "Item85  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent85 , golden_yjp85 , dut_yjp85 );
$fwrite(tri_report_ieee754, "Item86  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent86 , golden_yjp86 , dut_yjp86 );
$fwrite(tri_report_ieee754, "Item87  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent87 , golden_yjp87 , dut_yjp87 );
$fwrite(tri_report_ieee754, "Item88  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent88 , golden_yjp88 , dut_yjp88 );
$fwrite(tri_report_ieee754, "Item89  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent89 , golden_yjp89 , dut_yjp89 );
$fwrite(tri_report_ieee754, "Item90  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent90 , golden_yjp90 , dut_yjp90 );
$fwrite(tri_report_ieee754, "Item91  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent91 , golden_yjp91 , dut_yjp91 );
$fwrite(tri_report_ieee754, "Item92  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent92 , golden_yjp92 , dut_yjp92 );
$fwrite(tri_report_ieee754, "Item93  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent93 , golden_yjp93 , dut_yjp93 );
$fwrite(tri_report_ieee754, "Item94  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent94 , golden_yjp94 , dut_yjp94 );
$fwrite(tri_report_ieee754, "Item95  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent95 , golden_yjp95 , dut_yjp95 );
$fwrite(tri_report_ieee754, "Item96  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent96 , golden_yjp96 , dut_yjp96 );
$fwrite(tri_report_ieee754, "Item97  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent97 , golden_yjp97 , dut_yjp97 );
$fwrite(tri_report_ieee754, "Item98  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent98 , golden_yjp98 , dut_yjp98 );
$fwrite(tri_report_ieee754, "Item99  error percent: %f%%, golden result: %h, dut result: %h\n", error_percent99 , golden_yjp99 , dut_yjp99 );
$fwrite(tri_report_ieee754, "Item100 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent100, golden_yjp100, dut_yjp100);
$fwrite(tri_report_ieee754, "Item101 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent101, golden_yjp101, dut_yjp101);
$fwrite(tri_report_ieee754, "Item102 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent102, golden_yjp102, dut_yjp102);
$fwrite(tri_report_ieee754, "Item103 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent103, golden_yjp103, dut_yjp103);
$fwrite(tri_report_ieee754, "Item104 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent104, golden_yjp104, dut_yjp104);
$fwrite(tri_report_ieee754, "Item105 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent105, golden_yjp105, dut_yjp105);
$fwrite(tri_report_ieee754, "Item106 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent106, golden_yjp106, dut_yjp106);
$fwrite(tri_report_ieee754, "Item107 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent107, golden_yjp107, dut_yjp107);
$fwrite(tri_report_ieee754, "Item108 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent108, golden_yjp108, dut_yjp108);
$fwrite(tri_report_ieee754, "Item109 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent109, golden_yjp109, dut_yjp109);
$fwrite(tri_report_ieee754, "Item110 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent110, golden_yjp110, dut_yjp110);
$fwrite(tri_report_ieee754, "Item111 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent111, golden_yjp111, dut_yjp111);
$fwrite(tri_report_ieee754, "Item112 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent112, golden_yjp112, dut_yjp112);
$fwrite(tri_report_ieee754, "Item113 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent113, golden_yjp113, dut_yjp113);
$fwrite(tri_report_ieee754, "Item114 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent114, golden_yjp114, dut_yjp114);
$fwrite(tri_report_ieee754, "Item115 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent115, golden_yjp115, dut_yjp115);
$fwrite(tri_report_ieee754, "Item116 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent116, golden_yjp116, dut_yjp116);
$fwrite(tri_report_ieee754, "Item117 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent117, golden_yjp117, dut_yjp117);
$fwrite(tri_report_ieee754, "Item118 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent118, golden_yjp118, dut_yjp118);
$fwrite(tri_report_ieee754, "Item119 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent119, golden_yjp119, dut_yjp119);
$fwrite(tri_report_ieee754, "Item120 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent120, golden_yjp120, dut_yjp120);
$fwrite(tri_report_ieee754, "Item121 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent121, golden_yjp121, dut_yjp121);
$fwrite(tri_report_ieee754, "Item122 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent122, golden_yjp122, dut_yjp122);
$fwrite(tri_report_ieee754, "Item123 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent123, golden_yjp123, dut_yjp123);
$fwrite(tri_report_ieee754, "Item124 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent124, golden_yjp124, dut_yjp124);
$fwrite(tri_report_ieee754, "Item125 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent125, golden_yjp125, dut_yjp125);
$fwrite(tri_report_ieee754, "Item126 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent126, golden_yjp126, dut_yjp126);
$fwrite(tri_report_ieee754, "Item127 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent127, golden_yjp127, dut_yjp127);
$fwrite(tri_report_ieee754, "Item127 error percent: %f%%, golden result: %h, dut result: %h\n", error_percent127, golden_yjp127, dut_yjp127);
`endif //ST_WIDTH_INF_256
