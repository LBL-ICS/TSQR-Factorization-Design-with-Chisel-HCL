`ifdef ST_WIDTH_INF_16
$fwrite(tri_report, "===============================%d Column Results    ======================================\n",col_index);
if(col_index>=0  ) begin if(error_percent0  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item0   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent0  , ieee754_to_fp(golden_yjp0  ), ieee754_to_fp(dut_yjp0  )); end else begin $fwrite(tri_report, "Item0   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent0  , ieee754_to_fp(golden_yjp0  ), ieee754_to_fp(dut_yjp0  )); end end
if(col_index>=1  ) begin if(error_percent1  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item1   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent1  , ieee754_to_fp(golden_yjp1  ), ieee754_to_fp(dut_yjp1  )); end else begin $fwrite(tri_report, "Item1   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent1  , ieee754_to_fp(golden_yjp1  ), ieee754_to_fp(dut_yjp1  )); end end
if(col_index>=2  ) begin if(error_percent2  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item2   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent2  , ieee754_to_fp(golden_yjp2  ), ieee754_to_fp(dut_yjp2  )); end else begin $fwrite(tri_report, "Item2   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent2  , ieee754_to_fp(golden_yjp2  ), ieee754_to_fp(dut_yjp2  )); end end
if(col_index>=3  ) begin if(error_percent3  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item3   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent3  , ieee754_to_fp(golden_yjp3  ), ieee754_to_fp(dut_yjp3  )); end else begin $fwrite(tri_report, "Item3   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent3  , ieee754_to_fp(golden_yjp3  ), ieee754_to_fp(dut_yjp3  )); end end
if(col_index>=4  ) begin if(error_percent4  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item4   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent4  , ieee754_to_fp(golden_yjp4  ), ieee754_to_fp(dut_yjp4  )); end else begin $fwrite(tri_report, "Item4   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent4  , ieee754_to_fp(golden_yjp4  ), ieee754_to_fp(dut_yjp4  )); end end
if(col_index>=5  ) begin if(error_percent5  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item5   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent5  , ieee754_to_fp(golden_yjp5  ), ieee754_to_fp(dut_yjp5  )); end else begin $fwrite(tri_report, "Item5   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent5  , ieee754_to_fp(golden_yjp5  ), ieee754_to_fp(dut_yjp5  )); end end
if(col_index>=6  ) begin if(error_percent6  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item6   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent6  , ieee754_to_fp(golden_yjp6  ), ieee754_to_fp(dut_yjp6  )); end else begin $fwrite(tri_report, "Item6   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent6  , ieee754_to_fp(golden_yjp6  ), ieee754_to_fp(dut_yjp6  )); end end
if(col_index>=7  ) begin if(error_percent7  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item7   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent7  , ieee754_to_fp(golden_yjp7  ), ieee754_to_fp(dut_yjp7  )); end else begin $fwrite(tri_report, "Item7   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent7  , ieee754_to_fp(golden_yjp7  ), ieee754_to_fp(dut_yjp7  )); end end
`endif // ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32
if(col_index>=8  ) begin if(error_percent8  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item8   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent8  , ieee754_to_fp(golden_yjp8  ), ieee754_to_fp(dut_yjp8  )); end else begin $fwrite(tri_report, "Item8   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent8  , ieee754_to_fp(golden_yjp8  ), ieee754_to_fp(dut_yjp8  )); end end
if(col_index>=9  ) begin if(error_percent9  <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item9   Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent9  , ieee754_to_fp(golden_yjp9  ), ieee754_to_fp(dut_yjp9  )); end else begin $fwrite(tri_report, "Item9   Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent9  , ieee754_to_fp(golden_yjp9  ), ieee754_to_fp(dut_yjp9  )); end end
if(col_index>=10 ) begin if(error_percent10 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item10  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent10 , ieee754_to_fp(golden_yjp10 ), ieee754_to_fp(dut_yjp10 )); end else begin $fwrite(tri_report, "Item10  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent10 , ieee754_to_fp(golden_yjp10 ), ieee754_to_fp(dut_yjp10 )); end end
if(col_index>=11 ) begin if(error_percent11 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item11  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent11 , ieee754_to_fp(golden_yjp11 ), ieee754_to_fp(dut_yjp11 )); end else begin $fwrite(tri_report, "Item11  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent11 , ieee754_to_fp(golden_yjp11 ), ieee754_to_fp(dut_yjp11 )); end end
if(col_index>=12 ) begin if(error_percent12 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item12  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent12 , ieee754_to_fp(golden_yjp12 ), ieee754_to_fp(dut_yjp12 )); end else begin $fwrite(tri_report, "Item12  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent12 , ieee754_to_fp(golden_yjp12 ), ieee754_to_fp(dut_yjp12 )); end end
if(col_index>=13 ) begin if(error_percent13 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item13  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent13 , ieee754_to_fp(golden_yjp13 ), ieee754_to_fp(dut_yjp13 )); end else begin $fwrite(tri_report, "Item13  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent13 , ieee754_to_fp(golden_yjp13 ), ieee754_to_fp(dut_yjp13 )); end end
if(col_index>=14 ) begin if(error_percent14 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item14  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent14 , ieee754_to_fp(golden_yjp14 ), ieee754_to_fp(dut_yjp14 )); end else begin $fwrite(tri_report, "Item14  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent14 , ieee754_to_fp(golden_yjp14 ), ieee754_to_fp(dut_yjp14 )); end end
if(col_index>=15 ) begin if(error_percent15 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item15  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent15 , ieee754_to_fp(golden_yjp15 ), ieee754_to_fp(dut_yjp15 )); end else begin $fwrite(tri_report, "Item15  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent15 , ieee754_to_fp(golden_yjp15 ), ieee754_to_fp(dut_yjp15 )); end end
`endif // ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64
if(col_index>=16 ) begin if(error_percent16 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item16  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent16 , ieee754_to_fp(golden_yjp16 ), ieee754_to_fp(dut_yjp16 )); end else begin $fwrite(tri_report, "Item16  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent16 , ieee754_to_fp(golden_yjp16 ), ieee754_to_fp(dut_yjp16 )); end end
if(col_index>=17 ) begin if(error_percent17 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item17  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent17 , ieee754_to_fp(golden_yjp17 ), ieee754_to_fp(dut_yjp17 )); end else begin $fwrite(tri_report, "Item17  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent17 , ieee754_to_fp(golden_yjp17 ), ieee754_to_fp(dut_yjp17 )); end end
if(col_index>=18 ) begin if(error_percent18 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item18  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent18 , ieee754_to_fp(golden_yjp18 ), ieee754_to_fp(dut_yjp18 )); end else begin $fwrite(tri_report, "Item18  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent18 , ieee754_to_fp(golden_yjp18 ), ieee754_to_fp(dut_yjp18 )); end end
if(col_index>=19 ) begin if(error_percent19 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item19  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent19 , ieee754_to_fp(golden_yjp19 ), ieee754_to_fp(dut_yjp19 )); end else begin $fwrite(tri_report, "Item19  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent19 , ieee754_to_fp(golden_yjp19 ), ieee754_to_fp(dut_yjp19 )); end end
if(col_index>=20 ) begin if(error_percent20 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item20  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent20 , ieee754_to_fp(golden_yjp20 ), ieee754_to_fp(dut_yjp20 )); end else begin $fwrite(tri_report, "Item20  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent20 , ieee754_to_fp(golden_yjp20 ), ieee754_to_fp(dut_yjp20 )); end end
if(col_index>=21 ) begin if(error_percent21 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item21  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent21 , ieee754_to_fp(golden_yjp21 ), ieee754_to_fp(dut_yjp21 )); end else begin $fwrite(tri_report, "Item21  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent21 , ieee754_to_fp(golden_yjp21 ), ieee754_to_fp(dut_yjp21 )); end end
if(col_index>=22 ) begin if(error_percent22 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item22  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent22 , ieee754_to_fp(golden_yjp22 ), ieee754_to_fp(dut_yjp22 )); end else begin $fwrite(tri_report, "Item22  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent22 , ieee754_to_fp(golden_yjp22 ), ieee754_to_fp(dut_yjp22 )); end end
if(col_index>=23 ) begin if(error_percent23 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item23  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent23 , ieee754_to_fp(golden_yjp23 ), ieee754_to_fp(dut_yjp23 )); end else begin $fwrite(tri_report, "Item23  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent23 , ieee754_to_fp(golden_yjp23 ), ieee754_to_fp(dut_yjp23 )); end end
if(col_index>=24 ) begin if(error_percent24 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item24  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent24 , ieee754_to_fp(golden_yjp24 ), ieee754_to_fp(dut_yjp24 )); end else begin $fwrite(tri_report, "Item24  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent24 , ieee754_to_fp(golden_yjp24 ), ieee754_to_fp(dut_yjp24 )); end end
if(col_index>=25 ) begin if(error_percent25 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item25  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent25 , ieee754_to_fp(golden_yjp25 ), ieee754_to_fp(dut_yjp25 )); end else begin $fwrite(tri_report, "Item25  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent25 , ieee754_to_fp(golden_yjp25 ), ieee754_to_fp(dut_yjp25 )); end end
if(col_index>=26 ) begin if(error_percent26 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item26  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent26 , ieee754_to_fp(golden_yjp26 ), ieee754_to_fp(dut_yjp26 )); end else begin $fwrite(tri_report, "Item26  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent26 , ieee754_to_fp(golden_yjp26 ), ieee754_to_fp(dut_yjp26 )); end end
if(col_index>=27 ) begin if(error_percent27 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item27  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent27 , ieee754_to_fp(golden_yjp27 ), ieee754_to_fp(dut_yjp27 )); end else begin $fwrite(tri_report, "Item27  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent27 , ieee754_to_fp(golden_yjp27 ), ieee754_to_fp(dut_yjp27 )); end end
if(col_index>=28 ) begin if(error_percent28 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item28  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent28 , ieee754_to_fp(golden_yjp28 ), ieee754_to_fp(dut_yjp28 )); end else begin $fwrite(tri_report, "Item28  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent28 , ieee754_to_fp(golden_yjp28 ), ieee754_to_fp(dut_yjp28 )); end end
if(col_index>=29 ) begin if(error_percent29 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item29  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent29 , ieee754_to_fp(golden_yjp29 ), ieee754_to_fp(dut_yjp29 )); end else begin $fwrite(tri_report, "Item29  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent29 , ieee754_to_fp(golden_yjp29 ), ieee754_to_fp(dut_yjp29 )); end end
if(col_index>=30 ) begin if(error_percent30 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item30  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent30 , ieee754_to_fp(golden_yjp30 ), ieee754_to_fp(dut_yjp30 )); end else begin $fwrite(tri_report, "Item30  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent30 , ieee754_to_fp(golden_yjp30 ), ieee754_to_fp(dut_yjp30 )); end end
if(col_index>=31 ) begin if(error_percent31 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item31  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent31 , ieee754_to_fp(golden_yjp31 ), ieee754_to_fp(dut_yjp31 )); end else begin $fwrite(tri_report, "Item31  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent31 , ieee754_to_fp(golden_yjp31 ), ieee754_to_fp(dut_yjp31 )); end end
`endif // ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128
if(col_index>=32 ) begin if(error_percent32 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item32  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent32 , ieee754_to_fp(golden_yjp32 ), ieee754_to_fp(dut_yjp32 )); end else begin $fwrite(tri_report, "Item32  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent32 , ieee754_to_fp(golden_yjp32 ), ieee754_to_fp(dut_yjp32 )); end end
if(col_index>=33 ) begin if(error_percent33 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item33  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent33 , ieee754_to_fp(golden_yjp33 ), ieee754_to_fp(dut_yjp33 )); end else begin $fwrite(tri_report, "Item33  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent33 , ieee754_to_fp(golden_yjp33 ), ieee754_to_fp(dut_yjp33 )); end end
if(col_index>=34 ) begin if(error_percent34 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item34  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent34 , ieee754_to_fp(golden_yjp34 ), ieee754_to_fp(dut_yjp34 )); end else begin $fwrite(tri_report, "Item34  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent34 , ieee754_to_fp(golden_yjp34 ), ieee754_to_fp(dut_yjp34 )); end end
if(col_index>=35 ) begin if(error_percent35 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item35  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent35 , ieee754_to_fp(golden_yjp35 ), ieee754_to_fp(dut_yjp35 )); end else begin $fwrite(tri_report, "Item35  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent35 , ieee754_to_fp(golden_yjp35 ), ieee754_to_fp(dut_yjp35 )); end end
if(col_index>=36 ) begin if(error_percent36 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item36  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent36 , ieee754_to_fp(golden_yjp36 ), ieee754_to_fp(dut_yjp36 )); end else begin $fwrite(tri_report, "Item36  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent36 , ieee754_to_fp(golden_yjp36 ), ieee754_to_fp(dut_yjp36 )); end end
if(col_index>=37 ) begin if(error_percent37 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item37  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent37 , ieee754_to_fp(golden_yjp37 ), ieee754_to_fp(dut_yjp37 )); end else begin $fwrite(tri_report, "Item37  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent37 , ieee754_to_fp(golden_yjp37 ), ieee754_to_fp(dut_yjp37 )); end end
if(col_index>=38 ) begin if(error_percent38 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item38  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent38 , ieee754_to_fp(golden_yjp38 ), ieee754_to_fp(dut_yjp38 )); end else begin $fwrite(tri_report, "Item38  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent38 , ieee754_to_fp(golden_yjp38 ), ieee754_to_fp(dut_yjp38 )); end end
if(col_index>=39 ) begin if(error_percent39 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item39  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent39 , ieee754_to_fp(golden_yjp39 ), ieee754_to_fp(dut_yjp39 )); end else begin $fwrite(tri_report, "Item39  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent39 , ieee754_to_fp(golden_yjp39 ), ieee754_to_fp(dut_yjp39 )); end end
if(col_index>=40 ) begin if(error_percent40 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item40  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent40 , ieee754_to_fp(golden_yjp40 ), ieee754_to_fp(dut_yjp40 )); end else begin $fwrite(tri_report, "Item40  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent40 , ieee754_to_fp(golden_yjp40 ), ieee754_to_fp(dut_yjp40 )); end end
if(col_index>=41 ) begin if(error_percent41 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item41  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent41 , ieee754_to_fp(golden_yjp41 ), ieee754_to_fp(dut_yjp41 )); end else begin $fwrite(tri_report, "Item41  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent41 , ieee754_to_fp(golden_yjp41 ), ieee754_to_fp(dut_yjp41 )); end end
if(col_index>=42 ) begin if(error_percent42 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item42  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent42 , ieee754_to_fp(golden_yjp42 ), ieee754_to_fp(dut_yjp42 )); end else begin $fwrite(tri_report, "Item42  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent42 , ieee754_to_fp(golden_yjp42 ), ieee754_to_fp(dut_yjp42 )); end end
if(col_index>=43 ) begin if(error_percent43 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item43  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent43 , ieee754_to_fp(golden_yjp43 ), ieee754_to_fp(dut_yjp43 )); end else begin $fwrite(tri_report, "Item43  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent43 , ieee754_to_fp(golden_yjp43 ), ieee754_to_fp(dut_yjp43 )); end end
if(col_index>=44 ) begin if(error_percent44 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item44  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent44 , ieee754_to_fp(golden_yjp44 ), ieee754_to_fp(dut_yjp44 )); end else begin $fwrite(tri_report, "Item44  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent44 , ieee754_to_fp(golden_yjp44 ), ieee754_to_fp(dut_yjp44 )); end end
if(col_index>=45 ) begin if(error_percent45 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item45  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent45 , ieee754_to_fp(golden_yjp45 ), ieee754_to_fp(dut_yjp45 )); end else begin $fwrite(tri_report, "Item45  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent45 , ieee754_to_fp(golden_yjp45 ), ieee754_to_fp(dut_yjp45 )); end end
if(col_index>=46 ) begin if(error_percent46 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item46  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent46 , ieee754_to_fp(golden_yjp46 ), ieee754_to_fp(dut_yjp46 )); end else begin $fwrite(tri_report, "Item46  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent46 , ieee754_to_fp(golden_yjp46 ), ieee754_to_fp(dut_yjp46 )); end end
if(col_index>=47 ) begin if(error_percent47 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item47  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent47 , ieee754_to_fp(golden_yjp47 ), ieee754_to_fp(dut_yjp47 )); end else begin $fwrite(tri_report, "Item47  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent47 , ieee754_to_fp(golden_yjp47 ), ieee754_to_fp(dut_yjp47 )); end end
if(col_index>=48 ) begin if(error_percent48 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item48  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent48 , ieee754_to_fp(golden_yjp48 ), ieee754_to_fp(dut_yjp48 )); end else begin $fwrite(tri_report, "Item48  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent48 , ieee754_to_fp(golden_yjp48 ), ieee754_to_fp(dut_yjp48 )); end end
if(col_index>=49 ) begin if(error_percent49 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item49  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent49 , ieee754_to_fp(golden_yjp49 ), ieee754_to_fp(dut_yjp49 )); end else begin $fwrite(tri_report, "Item49  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent49 , ieee754_to_fp(golden_yjp49 ), ieee754_to_fp(dut_yjp49 )); end end
if(col_index>=50 ) begin if(error_percent50 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item50  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent50 , ieee754_to_fp(golden_yjp50 ), ieee754_to_fp(dut_yjp50 )); end else begin $fwrite(tri_report, "Item50  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent50 , ieee754_to_fp(golden_yjp50 ), ieee754_to_fp(dut_yjp50 )); end end
if(col_index>=51 ) begin if(error_percent51 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item51  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent51 , ieee754_to_fp(golden_yjp51 ), ieee754_to_fp(dut_yjp51 )); end else begin $fwrite(tri_report, "Item51  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent51 , ieee754_to_fp(golden_yjp51 ), ieee754_to_fp(dut_yjp51 )); end end
if(col_index>=52 ) begin if(error_percent52 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item52  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent52 , ieee754_to_fp(golden_yjp52 ), ieee754_to_fp(dut_yjp52 )); end else begin $fwrite(tri_report, "Item52  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent52 , ieee754_to_fp(golden_yjp52 ), ieee754_to_fp(dut_yjp52 )); end end
if(col_index>=53 ) begin if(error_percent53 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item53  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent53 , ieee754_to_fp(golden_yjp53 ), ieee754_to_fp(dut_yjp53 )); end else begin $fwrite(tri_report, "Item53  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent53 , ieee754_to_fp(golden_yjp53 ), ieee754_to_fp(dut_yjp53 )); end end
if(col_index>=54 ) begin if(error_percent54 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item54  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent54 , ieee754_to_fp(golden_yjp54 ), ieee754_to_fp(dut_yjp54 )); end else begin $fwrite(tri_report, "Item54  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent54 , ieee754_to_fp(golden_yjp54 ), ieee754_to_fp(dut_yjp54 )); end end
if(col_index>=55 ) begin if(error_percent55 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item55  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent55 , ieee754_to_fp(golden_yjp55 ), ieee754_to_fp(dut_yjp55 )); end else begin $fwrite(tri_report, "Item55  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent55 , ieee754_to_fp(golden_yjp55 ), ieee754_to_fp(dut_yjp55 )); end end
if(col_index>=56 ) begin if(error_percent56 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item56  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent56 , ieee754_to_fp(golden_yjp56 ), ieee754_to_fp(dut_yjp56 )); end else begin $fwrite(tri_report, "Item56  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent56 , ieee754_to_fp(golden_yjp56 ), ieee754_to_fp(dut_yjp56 )); end end
if(col_index>=57 ) begin if(error_percent57 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item57  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent57 , ieee754_to_fp(golden_yjp57 ), ieee754_to_fp(dut_yjp57 )); end else begin $fwrite(tri_report, "Item57  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent57 , ieee754_to_fp(golden_yjp57 ), ieee754_to_fp(dut_yjp57 )); end end
if(col_index>=58 ) begin if(error_percent58 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item58  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent58 , ieee754_to_fp(golden_yjp58 ), ieee754_to_fp(dut_yjp58 )); end else begin $fwrite(tri_report, "Item58  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent58 , ieee754_to_fp(golden_yjp58 ), ieee754_to_fp(dut_yjp58 )); end end
if(col_index>=59 ) begin if(error_percent59 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item59  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent59 , ieee754_to_fp(golden_yjp59 ), ieee754_to_fp(dut_yjp59 )); end else begin $fwrite(tri_report, "Item59  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent59 , ieee754_to_fp(golden_yjp59 ), ieee754_to_fp(dut_yjp59 )); end end
if(col_index>=60 ) begin if(error_percent60 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item60  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent60 , ieee754_to_fp(golden_yjp60 ), ieee754_to_fp(dut_yjp60 )); end else begin $fwrite(tri_report, "Item60  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent60 , ieee754_to_fp(golden_yjp60 ), ieee754_to_fp(dut_yjp60 )); end end
if(col_index>=61 ) begin if(error_percent61 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item61  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent61 , ieee754_to_fp(golden_yjp61 ), ieee754_to_fp(dut_yjp61 )); end else begin $fwrite(tri_report, "Item61  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent61 , ieee754_to_fp(golden_yjp61 ), ieee754_to_fp(dut_yjp61 )); end end
if(col_index>=62 ) begin if(error_percent62 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item62  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent62 , ieee754_to_fp(golden_yjp62 ), ieee754_to_fp(dut_yjp62 )); end else begin $fwrite(tri_report, "Item62  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent62 , ieee754_to_fp(golden_yjp62 ), ieee754_to_fp(dut_yjp62 )); end end
if(col_index>=63 ) begin if(error_percent63 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item63  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent63 , ieee754_to_fp(golden_yjp63 ), ieee754_to_fp(dut_yjp63 )); end else begin $fwrite(tri_report, "Item63  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent63 , ieee754_to_fp(golden_yjp63 ), ieee754_to_fp(dut_yjp63 )); end end
`endif // ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256
if(col_index>=64 ) begin if(error_percent64 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item64  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent64 , ieee754_to_fp(golden_yjp64 ), ieee754_to_fp(dut_yjp64 )); end else begin $fwrite(tri_report, "Item64  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent64 , ieee754_to_fp(golden_yjp64 ), ieee754_to_fp(dut_yjp64 )); end end
if(col_index>=65 ) begin if(error_percent65 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item65  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent65 , ieee754_to_fp(golden_yjp65 ), ieee754_to_fp(dut_yjp65 )); end else begin $fwrite(tri_report, "Item65  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent65 , ieee754_to_fp(golden_yjp65 ), ieee754_to_fp(dut_yjp65 )); end end
if(col_index>=66 ) begin if(error_percent66 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item66  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent66 , ieee754_to_fp(golden_yjp66 ), ieee754_to_fp(dut_yjp66 )); end else begin $fwrite(tri_report, "Item66  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent66 , ieee754_to_fp(golden_yjp66 ), ieee754_to_fp(dut_yjp66 )); end end
if(col_index>=67 ) begin if(error_percent67 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item67  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent67 , ieee754_to_fp(golden_yjp67 ), ieee754_to_fp(dut_yjp67 )); end else begin $fwrite(tri_report, "Item67  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent67 , ieee754_to_fp(golden_yjp67 ), ieee754_to_fp(dut_yjp67 )); end end
if(col_index>=68 ) begin if(error_percent68 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item68  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent68 , ieee754_to_fp(golden_yjp68 ), ieee754_to_fp(dut_yjp68 )); end else begin $fwrite(tri_report, "Item68  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent68 , ieee754_to_fp(golden_yjp68 ), ieee754_to_fp(dut_yjp68 )); end end
if(col_index>=69 ) begin if(error_percent69 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item69  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent69 , ieee754_to_fp(golden_yjp69 ), ieee754_to_fp(dut_yjp69 )); end else begin $fwrite(tri_report, "Item69  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent69 , ieee754_to_fp(golden_yjp69 ), ieee754_to_fp(dut_yjp69 )); end end
if(col_index>=70 ) begin if(error_percent70 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item70  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent70 , ieee754_to_fp(golden_yjp70 ), ieee754_to_fp(dut_yjp70 )); end else begin $fwrite(tri_report, "Item70  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent70 , ieee754_to_fp(golden_yjp70 ), ieee754_to_fp(dut_yjp70 )); end end
if(col_index>=71 ) begin if(error_percent71 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item71  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent71 , ieee754_to_fp(golden_yjp71 ), ieee754_to_fp(dut_yjp71 )); end else begin $fwrite(tri_report, "Item71  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent71 , ieee754_to_fp(golden_yjp71 ), ieee754_to_fp(dut_yjp71 )); end end
if(col_index>=72 ) begin if(error_percent72 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item72  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent72 , ieee754_to_fp(golden_yjp72 ), ieee754_to_fp(dut_yjp72 )); end else begin $fwrite(tri_report, "Item72  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent72 , ieee754_to_fp(golden_yjp72 ), ieee754_to_fp(dut_yjp72 )); end end
if(col_index>=73 ) begin if(error_percent73 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item73  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent73 , ieee754_to_fp(golden_yjp73 ), ieee754_to_fp(dut_yjp73 )); end else begin $fwrite(tri_report, "Item73  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent73 , ieee754_to_fp(golden_yjp73 ), ieee754_to_fp(dut_yjp73 )); end end
if(col_index>=74 ) begin if(error_percent74 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item74  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent74 , ieee754_to_fp(golden_yjp74 ), ieee754_to_fp(dut_yjp74 )); end else begin $fwrite(tri_report, "Item74  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent74 , ieee754_to_fp(golden_yjp74 ), ieee754_to_fp(dut_yjp74 )); end end
if(col_index>=75 ) begin if(error_percent75 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item75  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent75 , ieee754_to_fp(golden_yjp75 ), ieee754_to_fp(dut_yjp75 )); end else begin $fwrite(tri_report, "Item75  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent75 , ieee754_to_fp(golden_yjp75 ), ieee754_to_fp(dut_yjp75 )); end end
if(col_index>=76 ) begin if(error_percent76 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item76  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent76 , ieee754_to_fp(golden_yjp76 ), ieee754_to_fp(dut_yjp76 )); end else begin $fwrite(tri_report, "Item76  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent76 , ieee754_to_fp(golden_yjp76 ), ieee754_to_fp(dut_yjp76 )); end end
if(col_index>=77 ) begin if(error_percent77 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item77  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent77 , ieee754_to_fp(golden_yjp77 ), ieee754_to_fp(dut_yjp77 )); end else begin $fwrite(tri_report, "Item77  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent77 , ieee754_to_fp(golden_yjp77 ), ieee754_to_fp(dut_yjp77 )); end end
if(col_index>=78 ) begin if(error_percent78 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item78  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent78 , ieee754_to_fp(golden_yjp78 ), ieee754_to_fp(dut_yjp78 )); end else begin $fwrite(tri_report, "Item78  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent78 , ieee754_to_fp(golden_yjp78 ), ieee754_to_fp(dut_yjp78 )); end end
if(col_index>=79 ) begin if(error_percent79 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item79  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent79 , ieee754_to_fp(golden_yjp79 ), ieee754_to_fp(dut_yjp79 )); end else begin $fwrite(tri_report, "Item79  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent79 , ieee754_to_fp(golden_yjp79 ), ieee754_to_fp(dut_yjp79 )); end end
if(col_index>=80 ) begin if(error_percent80 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item80  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent80 , ieee754_to_fp(golden_yjp80 ), ieee754_to_fp(dut_yjp80 )); end else begin $fwrite(tri_report, "Item80  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent80 , ieee754_to_fp(golden_yjp80 ), ieee754_to_fp(dut_yjp80 )); end end
if(col_index>=81 ) begin if(error_percent81 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item81  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent81 , ieee754_to_fp(golden_yjp81 ), ieee754_to_fp(dut_yjp81 )); end else begin $fwrite(tri_report, "Item81  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent81 , ieee754_to_fp(golden_yjp81 ), ieee754_to_fp(dut_yjp81 )); end end
if(col_index>=82 ) begin if(error_percent82 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item82  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent82 , ieee754_to_fp(golden_yjp82 ), ieee754_to_fp(dut_yjp82 )); end else begin $fwrite(tri_report, "Item82  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent82 , ieee754_to_fp(golden_yjp82 ), ieee754_to_fp(dut_yjp82 )); end end
if(col_index>=83 ) begin if(error_percent83 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item83  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent83 , ieee754_to_fp(golden_yjp83 ), ieee754_to_fp(dut_yjp83 )); end else begin $fwrite(tri_report, "Item83  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent83 , ieee754_to_fp(golden_yjp83 ), ieee754_to_fp(dut_yjp83 )); end end
if(col_index>=84 ) begin if(error_percent84 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item84  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent84 , ieee754_to_fp(golden_yjp84 ), ieee754_to_fp(dut_yjp84 )); end else begin $fwrite(tri_report, "Item84  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent84 , ieee754_to_fp(golden_yjp84 ), ieee754_to_fp(dut_yjp84 )); end end
if(col_index>=85 ) begin if(error_percent85 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item85  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent85 , ieee754_to_fp(golden_yjp85 ), ieee754_to_fp(dut_yjp85 )); end else begin $fwrite(tri_report, "Item85  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent85 , ieee754_to_fp(golden_yjp85 ), ieee754_to_fp(dut_yjp85 )); end end
if(col_index>=86 ) begin if(error_percent86 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item86  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent86 , ieee754_to_fp(golden_yjp86 ), ieee754_to_fp(dut_yjp86 )); end else begin $fwrite(tri_report, "Item86  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent86 , ieee754_to_fp(golden_yjp86 ), ieee754_to_fp(dut_yjp86 )); end end
if(col_index>=87 ) begin if(error_percent87 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item87  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent87 , ieee754_to_fp(golden_yjp87 ), ieee754_to_fp(dut_yjp87 )); end else begin $fwrite(tri_report, "Item87  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent87 , ieee754_to_fp(golden_yjp87 ), ieee754_to_fp(dut_yjp87 )); end end
if(col_index>=88 ) begin if(error_percent88 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item88  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent88 , ieee754_to_fp(golden_yjp88 ), ieee754_to_fp(dut_yjp88 )); end else begin $fwrite(tri_report, "Item88  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent88 , ieee754_to_fp(golden_yjp88 ), ieee754_to_fp(dut_yjp88 )); end end
if(col_index>=89 ) begin if(error_percent89 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item89  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent89 , ieee754_to_fp(golden_yjp89 ), ieee754_to_fp(dut_yjp89 )); end else begin $fwrite(tri_report, "Item89  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent89 , ieee754_to_fp(golden_yjp89 ), ieee754_to_fp(dut_yjp89 )); end end
if(col_index>=90 ) begin if(error_percent90 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item90  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent90 , ieee754_to_fp(golden_yjp90 ), ieee754_to_fp(dut_yjp90 )); end else begin $fwrite(tri_report, "Item90  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent90 , ieee754_to_fp(golden_yjp90 ), ieee754_to_fp(dut_yjp90 )); end end
if(col_index>=91 ) begin if(error_percent91 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item91  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent91 , ieee754_to_fp(golden_yjp91 ), ieee754_to_fp(dut_yjp91 )); end else begin $fwrite(tri_report, "Item91  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent91 , ieee754_to_fp(golden_yjp91 ), ieee754_to_fp(dut_yjp91 )); end end
if(col_index>=92 ) begin if(error_percent92 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item92  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent92 , ieee754_to_fp(golden_yjp92 ), ieee754_to_fp(dut_yjp92 )); end else begin $fwrite(tri_report, "Item92  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent92 , ieee754_to_fp(golden_yjp92 ), ieee754_to_fp(dut_yjp92 )); end end
if(col_index>=93 ) begin if(error_percent93 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item93  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent93 , ieee754_to_fp(golden_yjp93 ), ieee754_to_fp(dut_yjp93 )); end else begin $fwrite(tri_report, "Item93  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent93 , ieee754_to_fp(golden_yjp93 ), ieee754_to_fp(dut_yjp93 )); end end
if(col_index>=94 ) begin if(error_percent94 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item94  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent94 , ieee754_to_fp(golden_yjp94 ), ieee754_to_fp(dut_yjp94 )); end else begin $fwrite(tri_report, "Item94  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent94 , ieee754_to_fp(golden_yjp94 ), ieee754_to_fp(dut_yjp94 )); end end
if(col_index>=95 ) begin if(error_percent95 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item95  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent95 , ieee754_to_fp(golden_yjp95 ), ieee754_to_fp(dut_yjp95 )); end else begin $fwrite(tri_report, "Item95  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent95 , ieee754_to_fp(golden_yjp95 ), ieee754_to_fp(dut_yjp95 )); end end
if(col_index>=96 ) begin if(error_percent96 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item96  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent96 , ieee754_to_fp(golden_yjp96 ), ieee754_to_fp(dut_yjp96 )); end else begin $fwrite(tri_report, "Item96  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent96 , ieee754_to_fp(golden_yjp96 ), ieee754_to_fp(dut_yjp96 )); end end
if(col_index>=97 ) begin if(error_percent97 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item97  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent97 , ieee754_to_fp(golden_yjp97 ), ieee754_to_fp(dut_yjp97 )); end else begin $fwrite(tri_report, "Item97  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent97 , ieee754_to_fp(golden_yjp97 ), ieee754_to_fp(dut_yjp97 )); end end
if(col_index>=98 ) begin if(error_percent98 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item98  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent98 , ieee754_to_fp(golden_yjp98 ), ieee754_to_fp(dut_yjp98 )); end else begin $fwrite(tri_report, "Item98  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent98 , ieee754_to_fp(golden_yjp98 ), ieee754_to_fp(dut_yjp98 )); end end
if(col_index>=99 ) begin if(error_percent99 <=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item99  Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent99 , ieee754_to_fp(golden_yjp99 ), ieee754_to_fp(dut_yjp99 )); end else begin $fwrite(tri_report, "Item99  Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent99 , ieee754_to_fp(golden_yjp99 ), ieee754_to_fp(dut_yjp99 )); end end
if(col_index>=100) begin if(error_percent100<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item100 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent100, ieee754_to_fp(golden_yjp100), ieee754_to_fp(dut_yjp100)); end else begin $fwrite(tri_report, "Item100 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent100, ieee754_to_fp(golden_yjp100), ieee754_to_fp(dut_yjp100)); end end
if(col_index>=101) begin if(error_percent101<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item101 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent101, ieee754_to_fp(golden_yjp101), ieee754_to_fp(dut_yjp101)); end else begin $fwrite(tri_report, "Item101 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent101, ieee754_to_fp(golden_yjp101), ieee754_to_fp(dut_yjp101)); end end
if(col_index>=102) begin if(error_percent102<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item102 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent102, ieee754_to_fp(golden_yjp102), ieee754_to_fp(dut_yjp102)); end else begin $fwrite(tri_report, "Item102 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent102, ieee754_to_fp(golden_yjp102), ieee754_to_fp(dut_yjp102)); end end
if(col_index>=103) begin if(error_percent103<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item103 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent103, ieee754_to_fp(golden_yjp103), ieee754_to_fp(dut_yjp103)); end else begin $fwrite(tri_report, "Item103 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent103, ieee754_to_fp(golden_yjp103), ieee754_to_fp(dut_yjp103)); end end
if(col_index>=104) begin if(error_percent104<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item104 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent104, ieee754_to_fp(golden_yjp104), ieee754_to_fp(dut_yjp104)); end else begin $fwrite(tri_report, "Item104 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent104, ieee754_to_fp(golden_yjp104), ieee754_to_fp(dut_yjp104)); end end
if(col_index>=105) begin if(error_percent105<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item105 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent105, ieee754_to_fp(golden_yjp105), ieee754_to_fp(dut_yjp105)); end else begin $fwrite(tri_report, "Item105 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent105, ieee754_to_fp(golden_yjp105), ieee754_to_fp(dut_yjp105)); end end
if(col_index>=106) begin if(error_percent106<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item106 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent106, ieee754_to_fp(golden_yjp106), ieee754_to_fp(dut_yjp106)); end else begin $fwrite(tri_report, "Item106 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent106, ieee754_to_fp(golden_yjp106), ieee754_to_fp(dut_yjp106)); end end
if(col_index>=107) begin if(error_percent107<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item107 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent107, ieee754_to_fp(golden_yjp107), ieee754_to_fp(dut_yjp107)); end else begin $fwrite(tri_report, "Item107 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent107, ieee754_to_fp(golden_yjp107), ieee754_to_fp(dut_yjp107)); end end
if(col_index>=108) begin if(error_percent108<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item108 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent108, ieee754_to_fp(golden_yjp108), ieee754_to_fp(dut_yjp108)); end else begin $fwrite(tri_report, "Item108 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent108, ieee754_to_fp(golden_yjp108), ieee754_to_fp(dut_yjp108)); end end
if(col_index>=109) begin if(error_percent109<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item109 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent109, ieee754_to_fp(golden_yjp109), ieee754_to_fp(dut_yjp109)); end else begin $fwrite(tri_report, "Item109 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent109, ieee754_to_fp(golden_yjp109), ieee754_to_fp(dut_yjp109)); end end
if(col_index>=110) begin if(error_percent110<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item110 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent110, ieee754_to_fp(golden_yjp110), ieee754_to_fp(dut_yjp110)); end else begin $fwrite(tri_report, "Item110 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent110, ieee754_to_fp(golden_yjp110), ieee754_to_fp(dut_yjp110)); end end
if(col_index>=111) begin if(error_percent111<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item111 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent111, ieee754_to_fp(golden_yjp111), ieee754_to_fp(dut_yjp111)); end else begin $fwrite(tri_report, "Item111 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent111, ieee754_to_fp(golden_yjp111), ieee754_to_fp(dut_yjp111)); end end
if(col_index>=112) begin if(error_percent112<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item112 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent112, ieee754_to_fp(golden_yjp112), ieee754_to_fp(dut_yjp112)); end else begin $fwrite(tri_report, "Item112 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent112, ieee754_to_fp(golden_yjp112), ieee754_to_fp(dut_yjp112)); end end
if(col_index>=113) begin if(error_percent113<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item113 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent113, ieee754_to_fp(golden_yjp113), ieee754_to_fp(dut_yjp113)); end else begin $fwrite(tri_report, "Item113 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent113, ieee754_to_fp(golden_yjp113), ieee754_to_fp(dut_yjp113)); end end
if(col_index>=114) begin if(error_percent114<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item114 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent114, ieee754_to_fp(golden_yjp114), ieee754_to_fp(dut_yjp114)); end else begin $fwrite(tri_report, "Item114 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent114, ieee754_to_fp(golden_yjp114), ieee754_to_fp(dut_yjp114)); end end
if(col_index>=115) begin if(error_percent115<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item115 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent115, ieee754_to_fp(golden_yjp115), ieee754_to_fp(dut_yjp115)); end else begin $fwrite(tri_report, "Item115 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent115, ieee754_to_fp(golden_yjp115), ieee754_to_fp(dut_yjp115)); end end
if(col_index>=116) begin if(error_percent116<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item116 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent116, ieee754_to_fp(golden_yjp116), ieee754_to_fp(dut_yjp116)); end else begin $fwrite(tri_report, "Item116 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent116, ieee754_to_fp(golden_yjp116), ieee754_to_fp(dut_yjp116)); end end
if(col_index>=117) begin if(error_percent117<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item117 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent117, ieee754_to_fp(golden_yjp117), ieee754_to_fp(dut_yjp117)); end else begin $fwrite(tri_report, "Item117 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent117, ieee754_to_fp(golden_yjp117), ieee754_to_fp(dut_yjp117)); end end
if(col_index>=118) begin if(error_percent118<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item118 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent118, ieee754_to_fp(golden_yjp118), ieee754_to_fp(dut_yjp118)); end else begin $fwrite(tri_report, "Item118 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent118, ieee754_to_fp(golden_yjp118), ieee754_to_fp(dut_yjp118)); end end
if(col_index>=119) begin if(error_percent119<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item119 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent119, ieee754_to_fp(golden_yjp119), ieee754_to_fp(dut_yjp119)); end else begin $fwrite(tri_report, "Item119 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent119, ieee754_to_fp(golden_yjp119), ieee754_to_fp(dut_yjp119)); end end
if(col_index>=120) begin if(error_percent120<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item120 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent120, ieee754_to_fp(golden_yjp120), ieee754_to_fp(dut_yjp120)); end else begin $fwrite(tri_report, "Item120 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent120, ieee754_to_fp(golden_yjp120), ieee754_to_fp(dut_yjp120)); end end
if(col_index>=121) begin if(error_percent121<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item121 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent121, ieee754_to_fp(golden_yjp121), ieee754_to_fp(dut_yjp121)); end else begin $fwrite(tri_report, "Item121 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent121, ieee754_to_fp(golden_yjp121), ieee754_to_fp(dut_yjp121)); end end
if(col_index>=122) begin if(error_percent122<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item122 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent122, ieee754_to_fp(golden_yjp122), ieee754_to_fp(dut_yjp122)); end else begin $fwrite(tri_report, "Item122 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent122, ieee754_to_fp(golden_yjp122), ieee754_to_fp(dut_yjp122)); end end
if(col_index>=123) begin if(error_percent123<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item123 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent123, ieee754_to_fp(golden_yjp123), ieee754_to_fp(dut_yjp123)); end else begin $fwrite(tri_report, "Item123 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent123, ieee754_to_fp(golden_yjp123), ieee754_to_fp(dut_yjp123)); end end
if(col_index>=124) begin if(error_percent124<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item124 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent124, ieee754_to_fp(golden_yjp124), ieee754_to_fp(dut_yjp124)); end else begin $fwrite(tri_report, "Item124 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent124, ieee754_to_fp(golden_yjp124), ieee754_to_fp(dut_yjp124)); end end
if(col_index>=125) begin if(error_percent125<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item125 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent125, ieee754_to_fp(golden_yjp125), ieee754_to_fp(dut_yjp125)); end else begin $fwrite(tri_report, "Item125 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent125, ieee754_to_fp(golden_yjp125), ieee754_to_fp(dut_yjp125)); end end
if(col_index>=126) begin if(error_percent126<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item126 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent126, ieee754_to_fp(golden_yjp126), ieee754_to_fp(dut_yjp126)); end else begin $fwrite(tri_report, "Item126 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent126, ieee754_to_fp(golden_yjp126), ieee754_to_fp(dut_yjp126)); end end
if(col_index==127) begin if(error_percent127<=`ERROR_THRESHOLD) begin $fwrite(tri_report, "Item127 Comp Pass! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent127, ieee754_to_fp(golden_yjp127), ieee754_to_fp(dut_yjp127)); end else begin $fwrite(tri_report, "Item127 Comp FAIL! error percent: %f%%, golden result: %f, dut result: %f\n", error_percent127, ieee754_to_fp(golden_yjp127), ieee754_to_fp(dut_yjp127)); end end
`endif // ST_WIDTH_INF_256
