module fsm(
  input          clk,
  input          rst,
  input          tsqr_en,
  input  [15:0]  tile_no,
  output [15:0]  hh_cnt,
  output [15:0]  mx_cnt,
  output         d1_rdy,
  output         d1_vld,
  output         d2_vld,
  output         vk1_vld,
  output         d3_rdy,
  output         d3_vld,
  output         tk_vld,
  output         d4_rdy,
  output         d5_rdy,
  output         d5_vld,
  output         yj_sft,
  output         d4_sft,
  output         hh_st,
  output         mem0_fi,
  output         mem1_fi,
  output         tsqr_fi,
  output         dmx0_mem_ena,
  output [127:0] dmx0_mem_wea,
  output [4:0]   dmx0_mem_addra,
  output         dmx0_mem_enb,
  output [4:0]   dmx0_mem_addrb,
  output         dmx1_mem_ena,
  output [127:0] dmx1_mem_wea,
  output [4:0]   dmx1_mem_addra,
  output         dmx1_mem_enb,
  output [4:0]   dmx1_mem_addrb,
  output         rtri_mem_ena,
  output [127:0] rtri_mem_wea,
  output [4:0]   rtri_mem_addra,
  output         rtri_mem_enb,
  output [4:0]   rtri_mem_addrb
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [127:0] _RAND_23;
  reg [127:0] _RAND_24;
  reg [127:0] _RAND_25;
  reg [127:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
`endif // RANDOMIZE_REG_INIT
  reg  hh_en; // @[tsqr_fsm.scala 94:24]
  wire  _T = mem0_fi | mem1_fi; // @[tsqr_fsm.scala 98:28]
  wire  _GEN_0 = tsqr_en | hh_en; // @[tsqr_fsm.scala 100:28 101:19 94:24]
  reg [15:0] cnt; // @[tsqr_fsm.scala 104:22]
  reg [15:0] nxt_hh_cnt; // @[tsqr_fsm.scala 106:29]
  reg [15:0] nxt_mx_cnt; // @[tsqr_fsm.scala 107:29]
  wire  _T_1 = cnt == 16'h1f1; // @[tsqr_fsm.scala 109:18]
  wire [15:0] _nxt_cnt_T_1 = cnt + 16'h1; // @[tsqr_fsm.scala 112:28]
  wire [6:0] _T_3 = 7'h40 / 2'h2; // @[tsqr_fsm.scala 117:64]
  wire [6:0] _T_5 = _T_3 - 7'h1; // @[tsqr_fsm.scala 117:68]
  wire [15:0] _GEN_72 = {{9'd0}, _T_5}; // @[tsqr_fsm.scala 117:42]
  wire [15:0] _nxt_hh_cnt_T_1 = hh_cnt + 16'h1; // @[tsqr_fsm.scala 120:34]
  wire  _T_10 = hh_cnt == 16'h1f; // @[tsqr_fsm.scala 125:22]
  wire [15:0] _T_12 = tile_no - 16'h1; // @[tsqr_fsm.scala 125:72]
  wire  _T_13 = mx_cnt == _T_12; // @[tsqr_fsm.scala 125:59]
  wire [15:0] _nxt_mx_cnt_T_1 = mx_cnt + 16'h1; // @[tsqr_fsm.scala 128:34]
  reg [15:0] tr_cy_reg; // @[tsqr_fsm.scala 143:28]
  reg  tr_cnt_en; // @[tsqr_fsm.scala 144:28]
  reg [15:0] tr_cnt; // @[tsqr_fsm.scala 145:25]
  wire  rd_mem_fst = rst ? 1'h0 : tsqr_en & ~hh_en; // @[tsqr_fsm.scala 151:18 152:24 157:24]
  wire  wr_mem_st = rst ? 1'h0 : hh_en & tr_cnt == 16'hfa; // @[tsqr_fsm.scala 151:18 153:23 158:23]
  wire  rd_mem_st = rst ? 1'h0 : hh_en & cnt == 16'hf0; // @[tsqr_fsm.scala 151:18 155:23 160:23]
  wire [15:0] _tr_cy_T_1 = 16'h20 - hh_cnt; // @[tsqr_fsm.scala 166:45]
  wire [15:0] tr_cy = rd_mem_st ? _tr_cy_T_1 : tr_cy_reg; // @[tsqr_fsm.scala 165:24 166:19 168:19]
  wire [15:0] _hh_fi_T_1 = 16'hfb + tr_cy; // @[tsqr_fsm.scala 172:45]
  wire [15:0] _hh_fi_T_3 = _hh_fi_T_1 + 16'h1; // @[tsqr_fsm.scala 172:53]
  wire  hh_fi = tr_cnt == _hh_fi_T_3; // @[tsqr_fsm.scala 172:26]
  wire [15:0] _nxt_tr_cnt_T_1 = tr_cnt + 16'h1; // @[tsqr_fsm.scala 178:34]
  wire  _GEN_21 = hh_en & cnt == 16'hf4 | tr_cnt_en; // @[tsqr_fsm.scala 195:51 196:23 144:28]
  reg  d1_rdy_REG; // @[tsqr_fsm.scala 200:26]
  reg  d1_vld_REG; // @[tsqr_fsm.scala 201:26]
  reg  d2_vld_REG; // @[tsqr_fsm.scala 203:26]
  wire  _vk1_vld_T = cnt == 16'hf3; // @[tsqr_fsm.scala 205:41]
  reg  vk1_vld_REG; // @[tsqr_fsm.scala 205:27]
  reg  d3_rdy_REG; // @[tsqr_fsm.scala 206:26]
  reg  d3_vld_REG; // @[tsqr_fsm.scala 207:26]
  reg  tk_vld_REG; // @[tsqr_fsm.scala 209:26]
  wire  _d4_vld_T_1 = tr_cnt_en & tr_cnt >= 16'h5a; // @[tsqr_fsm.scala 212:29]
  wire [15:0] _d4_vld_T_3 = 16'h5a + tr_cy; // @[tsqr_fsm.scala 212:78]
  wire [15:0] _d5_rdy_T_7 = _d4_vld_T_3 + 16'h80; // @[tsqr_fsm.scala 213:100]
  wire [15:0] _d5_vld_T_11 = _d5_rdy_T_7 + 16'ha; // @[tsqr_fsm.scala 214:127]
  wire  _yjp_vld_T_16 = tr_cnt >= 16'hfb; // @[tsqr_fsm.scala 216:112]
  wire [15:0] _d4_sft_T_5 = 16'hda + tr_cy; // @[tsqr_fsm.scala 218:90]
  wire [15:0] _yj_sft_T_1 = 16'he3 + tr_cy; // @[tsqr_fsm.scala 219:54]
  reg  dmx0_mem_enb_reg; // @[tsqr_fsm.scala 250:35]
  reg  dmx1_mem_enb_reg; // @[tsqr_fsm.scala 251:35]
  reg  rtri_mem_enb_reg; // @[tsqr_fsm.scala 252:35]
  reg  dmx0_mem_ena_reg; // @[tsqr_fsm.scala 253:35]
  reg  dmx1_mem_ena_reg; // @[tsqr_fsm.scala 254:35]
  reg  rtri_mem_ena_reg; // @[tsqr_fsm.scala 255:35]
  wire  _rd_dmx0_en_T_1 = ~mx_cnt[0]; // @[tsqr_fsm.scala 269:27]
  wire [15:0] _rd_dmx0_en_T_4 = 16'hf2 + tr_cy; // @[tsqr_fsm.scala 269:76]
  wire  _rd_dmx0_en_T_6 = cnt >= 16'hf2 & cnt < _rd_dmx0_en_T_4; // @[tsqr_fsm.scala 269:58]
  wire  rd_dmx0_en = rst ? 1'h0 : ~mx_cnt[0] & (cnt >= 16'hf2 & cnt < _rd_dmx0_en_T_4); // @[tsqr_fsm.scala 261:18 262:24 269:24]
  wire  rd_dmx1_en = rst ? 1'h0 : mx_cnt[0] & _rd_dmx0_en_T_6; // @[tsqr_fsm.scala 261:18 263:24 270:24]
  wire  rd_rtri_en = rst ? 1'h0 : _rd_dmx0_en_T_6; // @[tsqr_fsm.scala 261:18 264:24 271:24]
  reg [4:0] dmx0_mem_addrb_reg; // @[tsqr_fsm.scala 277:37]
  reg [4:0] dmx1_mem_addrb_reg; // @[tsqr_fsm.scala 278:37]
  reg [4:0] rtri_mem_addrb_reg; // @[tsqr_fsm.scala 279:37]
  wire  _T_26 = hh_en & cnt == 16'hf2; // @[tsqr_fsm.scala 294:40]
  wire [4:0] _dmx0_mem_addrb_wire_T_1 = dmx0_mem_addrb_reg + 5'h1; // @[tsqr_fsm.scala 297:55]
  wire [4:0] _GEN_30 = rd_dmx0_en ? _dmx0_mem_addrb_wire_T_1 : dmx0_mem_addrb_reg; // @[tsqr_fsm.scala 296:31 297:33 299:33]
  wire [15:0] _GEN_31 = _rd_dmx0_en_T_1 & (hh_en & cnt == 16'hf2) ? hh_cnt : {{11'd0}, _GEN_30}; // @[tsqr_fsm.scala 294:63 295:32]
  wire [15:0] _GEN_32 = rd_mem_fst ? 16'h0 : _GEN_31; // @[tsqr_fsm.scala 292:25 293:33]
  wire [4:0] _dmx1_mem_addrb_wire_T_1 = dmx1_mem_addrb_reg + 5'h1; // @[tsqr_fsm.scala 307:55]
  wire [4:0] _GEN_33 = rd_dmx1_en ? _dmx1_mem_addrb_wire_T_1 : dmx1_mem_addrb_reg; // @[tsqr_fsm.scala 306:31 307:33 309:33]
  wire [15:0] _GEN_34 = mx_cnt[0] & _T_26 ? hh_cnt : {{11'd0}, _GEN_33}; // @[tsqr_fsm.scala 304:62 305:33]
  wire [15:0] _GEN_35 = rd_mem_fst ? 16'h0 : _GEN_34; // @[tsqr_fsm.scala 302:25 303:33]
  wire [4:0] _rtri_mem_addrb_wire_T_1 = rtri_mem_addrb_reg + 5'h1; // @[tsqr_fsm.scala 317:55]
  wire [4:0] _GEN_36 = rd_rtri_en ? _rtri_mem_addrb_wire_T_1 : rtri_mem_addrb_reg; // @[tsqr_fsm.scala 316:31 317:33 319:33]
  wire [15:0] _GEN_37 = _T_26 ? hh_cnt : {{11'd0}, _GEN_36}; // @[tsqr_fsm.scala 314:50 315:33]
  wire [15:0] _GEN_38 = rd_mem_fst ? 16'h0 : _GEN_37; // @[tsqr_fsm.scala 312:25 313:33]
  reg [127:0] dmx0_mem_wea_reg; // @[tsqr_fsm.scala 322:35]
  reg [127:0] dmx1_mem_wea_reg; // @[tsqr_fsm.scala 323:35]
  reg [127:0] rtri_mem_wea_reg; // @[tsqr_fsm.scala 324:35]
  reg [127:0] rtri_mem_wea_update; // @[tsqr_fsm.scala 327:38]
  wire  _dmx0_mem_ena_wire_T_6 = tr_cnt < _hh_fi_T_1; // @[tsqr_fsm.scala 334:85]
  wire  dmx0_mem_ena_wire = rst ? 1'h0 : _rd_dmx0_en_T_1 & _yjp_vld_T_16 & tr_cnt < _hh_fi_T_1; // @[tsqr_fsm.scala 329:18 330:31 334:31]
  wire  dmx1_mem_ena_wire = rst ? 1'h0 : mx_cnt[0] & _yjp_vld_T_16 & _dmx0_mem_ena_wire_T_6; // @[tsqr_fsm.scala 329:18 331:31 335:31]
  wire  rtri_mem_ena_wire = rst ? 1'h0 : _yjp_vld_T_16 & _dmx0_mem_ena_wire_T_6; // @[tsqr_fsm.scala 329:18 332:31 336:31]
  reg [4:0] dmx0_mem_addra_reg; // @[tsqr_fsm.scala 367:37]
  reg [4:0] dmx1_mem_addra_reg; // @[tsqr_fsm.scala 368:37]
  reg [4:0] rtri_mem_addra_reg; // @[tsqr_fsm.scala 369:37]
  wire  _T_42 = hh_en & tr_cnt == 16'hfb; // @[tsqr_fsm.scala 371:34]
  wire [4:0] _dmx0_mem_addra_wire_T_1 = dmx0_mem_addra_reg + 5'h1; // @[tsqr_fsm.scala 374:55]
  wire [4:0] _GEN_48 = dmx0_mem_ena_wire ? _dmx0_mem_addra_wire_T_1 : dmx0_mem_addra_reg; // @[tsqr_fsm.scala 373:38 374:33 376:33]
  wire [15:0] _GEN_49 = _rd_dmx0_en_T_1 & (hh_en & tr_cnt == 16'hfb) ? hh_cnt : {{11'd0}, _GEN_48}; // @[tsqr_fsm.scala 371:66 372:33]
  wire [4:0] _dmx1_mem_addra_wire_T_1 = dmx1_mem_addra_reg + 5'h1; // @[tsqr_fsm.scala 382:55]
  wire [4:0] _GEN_50 = dmx1_mem_ena_wire ? _dmx1_mem_addra_wire_T_1 : dmx1_mem_addra_reg; // @[tsqr_fsm.scala 381:38 382:33 384:33]
  wire [15:0] _GEN_51 = mx_cnt[0] & _T_42 ? hh_cnt : {{11'd0}, _GEN_50}; // @[tsqr_fsm.scala 379:65 380:33]
  wire [4:0] _rtri_mem_addra_wire_T_1 = rtri_mem_addra_reg + 5'h1; // @[tsqr_fsm.scala 390:55]
  wire [4:0] _GEN_52 = rtri_mem_ena_wire ? _rtri_mem_addra_wire_T_1 : rtri_mem_addra_reg; // @[tsqr_fsm.scala 389:38 390:33 392:33]
  wire [15:0] _GEN_53 = _T_42 ? hh_cnt : {{11'd0}, _GEN_52}; // @[tsqr_fsm.scala 387:53 388:33]
  wire [4:0] dmx0_mem_addra_wire = _GEN_49[4:0]; // @[tsqr_fsm.scala 286:39]
  wire [4:0] dmx1_mem_addra_wire = _GEN_51[4:0]; // @[tsqr_fsm.scala 287:39]
  wire [4:0] rtri_mem_addra_wire = _GEN_53[4:0]; // @[tsqr_fsm.scala 288:39]
  wire [4:0] dmx0_mem_addrb_wire = _GEN_32[4:0]; // @[tsqr_fsm.scala 283:39]
  wire [4:0] dmx1_mem_addrb_wire = _GEN_35[4:0]; // @[tsqr_fsm.scala 284:39]
  wire [4:0] rtri_mem_addrb_wire = _GEN_38[4:0]; // @[tsqr_fsm.scala 285:39]
  wire [16:0] _mem0_fi_T_4 = {{1'd0}, _hh_fi_T_1}; // @[tsqr_fsm.scala 435:63]
  wire  _mem0_fi_T_6 = tr_cnt == _mem0_fi_T_4[15:0]; // @[tsqr_fsm.scala 435:36]
  wire  _mem0_fi_T_8 = tr_cy == 16'h1; // @[tsqr_fsm.scala 435:80]
  wire [18:0] _rtri_mem_wea_update_T_2 = hh_cnt * 3'h4; // @[tsqr_fsm.scala 449:62]
  wire [127:0] _rtri_mem_wea_update_T_3 = rtri_mem_wea_update >> _rtri_mem_wea_update_T_2; // @[tsqr_fsm.scala 449:52]
  assign hh_cnt = rst ? 16'h0 : nxt_hh_cnt; // @[tsqr_fsm.scala 133:18 135:20 139:20]
  assign mx_cnt = rst ? 16'h0 : nxt_mx_cnt; // @[tsqr_fsm.scala 133:18 136:20 140:20]
  assign d1_rdy = d1_rdy_REG; // @[tsqr_fsm.scala 200:16]
  assign d1_vld = d1_vld_REG; // @[tsqr_fsm.scala 201:16]
  assign d2_vld = d2_vld_REG; // @[tsqr_fsm.scala 203:16]
  assign vk1_vld = vk1_vld_REG; // @[tsqr_fsm.scala 205:17]
  assign d3_rdy = d3_rdy_REG; // @[tsqr_fsm.scala 206:16]
  assign d3_vld = d3_vld_REG; // @[tsqr_fsm.scala 207:16]
  assign tk_vld = tk_vld_REG; // @[tsqr_fsm.scala 209:16]
  assign d4_rdy = tr_cnt_en & tr_cnt < tr_cy; // @[tsqr_fsm.scala 211:29]
  assign d5_rdy = tr_cnt_en & tr_cnt >= 16'hda & tr_cnt < _d5_rdy_T_7; // @[tsqr_fsm.scala 213:69]
  assign d5_vld = tr_cnt_en & tr_cnt >= 16'he4 & tr_cnt < _d5_vld_T_11; // @[tsqr_fsm.scala 214:82]
  assign yj_sft = tr_cnt_en & tr_cnt < _yj_sft_T_1; // @[tsqr_fsm.scala 219:28]
  assign d4_sft = _d4_vld_T_1 & tr_cnt < _d4_sft_T_5; // @[tsqr_fsm.scala 218:53]
  assign hh_st = rst ? 1'h0 : hh_en & tr_cnt == 16'hfd; // @[tsqr_fsm.scala 151:18 154:19 159:19]
  assign mem0_fi = _rd_dmx0_en_T_1 & tr_cnt == _mem0_fi_T_4[15:0] & tr_cy == 16'h1; // @[tsqr_fsm.scala 435:71]
  assign mem1_fi = mx_cnt[0] & _mem0_fi_T_6 & _mem0_fi_T_8; // @[tsqr_fsm.scala 436:69]
  assign tsqr_fi = _T & _T_13; // @[tsqr_fsm.scala 440:36]
  assign dmx0_mem_ena = dmx0_mem_ena_reg; // @[tsqr_fsm.scala 461:22]
  assign dmx0_mem_wea = _rd_dmx0_en_T_1 & wr_mem_st ? 128'hffffffffffffffffffffffffffffffff : dmx0_mem_wea_reg; // @[tsqr_fsm.scala 339:37 340:26 342:26]
  assign dmx0_mem_addra = dmx0_mem_addra_reg; // @[tsqr_fsm.scala 429:20]
  assign dmx0_mem_enb = dmx0_mem_enb_reg; // @[tsqr_fsm.scala 458:22]
  assign dmx0_mem_addrb = dmx0_mem_addrb_reg; // @[tsqr_fsm.scala 426:20]
  assign dmx1_mem_ena = dmx1_mem_ena_reg; // @[tsqr_fsm.scala 462:22]
  assign dmx1_mem_wea = mx_cnt[0] & wr_mem_st ? 128'hffffffffffffffffffffffffffffffff : dmx1_mem_wea_reg; // @[tsqr_fsm.scala 345:36 346:26 348:26]
  assign dmx1_mem_addra = dmx1_mem_addra_reg; // @[tsqr_fsm.scala 430:20]
  assign dmx1_mem_enb = dmx1_mem_enb_reg; // @[tsqr_fsm.scala 459:22]
  assign dmx1_mem_addrb = dmx1_mem_addrb_reg; // @[tsqr_fsm.scala 427:20]
  assign rtri_mem_ena = rtri_mem_ena_reg; // @[tsqr_fsm.scala 463:22]
  assign rtri_mem_wea = wr_mem_st ? rtri_mem_wea_update : rtri_mem_wea_reg; // @[tsqr_fsm.scala 351:24 352:26 354:26]
  assign rtri_mem_addra = rtri_mem_addra_reg; // @[tsqr_fsm.scala 431:20]
  assign rtri_mem_enb = rtri_mem_enb_reg; // @[tsqr_fsm.scala 460:22]
  assign rtri_mem_addrb = rtri_mem_addrb_reg; // @[tsqr_fsm.scala 428:20]
  always @(posedge clk) begin
    if (rst) begin // @[tsqr_fsm.scala 96:18]
      hh_en <= 1'h0; // @[tsqr_fsm.scala 97:19]
    end else if (mem0_fi | mem1_fi) begin // @[tsqr_fsm.scala 98:38]
      hh_en <= 1'h0; // @[tsqr_fsm.scala 99:19]
    end else begin
      hh_en <= _GEN_0;
    end
    if (rst) begin // @[tsqr_fsm.scala 133:18]
      cnt <= 16'h0; // @[tsqr_fsm.scala 134:17]
    end else if (cnt == 16'h1f1) begin // @[tsqr_fsm.scala 109:34]
      cnt <= 16'h0; // @[tsqr_fsm.scala 110:21]
    end else if (hh_en) begin // @[tsqr_fsm.scala 111:26]
      cnt <= _nxt_cnt_T_1; // @[tsqr_fsm.scala 112:21]
    end
    if (_T_1 & hh_cnt == _GEN_72) begin // @[tsqr_fsm.scala 117:75]
      nxt_hh_cnt <= 16'h0; // @[tsqr_fsm.scala 118:24]
    end else if (hh_en & _T_1) begin // @[tsqr_fsm.scala 119:48]
      nxt_hh_cnt <= _nxt_hh_cnt_T_1; // @[tsqr_fsm.scala 120:24]
    end else begin
      nxt_hh_cnt <= hh_cnt; // @[tsqr_fsm.scala 122:24]
    end
    if (hh_cnt == 16'h1f & mx_cnt == _T_12 & _T_1) begin // @[tsqr_fsm.scala 125:101]
      nxt_mx_cnt <= 16'h0; // @[tsqr_fsm.scala 126:24]
    end else if (hh_en & _T_10 & _T_1) begin // @[tsqr_fsm.scala 127:85]
      nxt_mx_cnt <= _nxt_mx_cnt_T_1; // @[tsqr_fsm.scala 128:24]
    end else begin
      nxt_mx_cnt <= mx_cnt; // @[tsqr_fsm.scala 130:24]
    end
    if (rst) begin // @[tsqr_fsm.scala 183:18]
      tr_cy_reg <= 16'h0; // @[tsqr_fsm.scala 185:23]
    end else if (rd_mem_st) begin // @[tsqr_fsm.scala 165:24]
      tr_cy_reg <= _tr_cy_T_1; // @[tsqr_fsm.scala 166:19]
    end
    if (rst) begin // @[tsqr_fsm.scala 191:18]
      tr_cnt_en <= 1'h0; // @[tsqr_fsm.scala 192:23]
    end else if (hh_fi) begin // @[tsqr_fsm.scala 193:26]
      tr_cnt_en <= 1'h0; // @[tsqr_fsm.scala 194:23]
    end else begin
      tr_cnt_en <= _GEN_21;
    end
    if (rst) begin // @[tsqr_fsm.scala 183:18]
      tr_cnt <= 16'h0; // @[tsqr_fsm.scala 184:20]
    end else if (hh_fi) begin // @[tsqr_fsm.scala 175:20]
      tr_cnt <= 16'h0; // @[tsqr_fsm.scala 176:24]
    end else if (tr_cnt_en) begin // @[tsqr_fsm.scala 177:30]
      tr_cnt <= _nxt_tr_cnt_T_1; // @[tsqr_fsm.scala 178:24]
    end
    d1_rdy_REG <= hh_en & cnt == 16'h1; // @[tsqr_fsm.scala 200:33]
    d1_vld_REG <= hh_en & cnt == 16'h5b; // @[tsqr_fsm.scala 201:33]
    d2_vld_REG <= hh_en & cnt == 16'he6; // @[tsqr_fsm.scala 203:33]
    vk1_vld_REG <= hh_en & cnt == 16'hf3; // @[tsqr_fsm.scala 205:34]
    d3_rdy_REG <= hh_en & _vk1_vld_T; // @[tsqr_fsm.scala 206:33]
    d3_vld_REG <= hh_en & cnt == 16'h14d; // @[tsqr_fsm.scala 207:33]
    tk_vld_REG <= hh_en & cnt == 16'h1ce; // @[tsqr_fsm.scala 209:33]
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx0_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 403:26]
    end else if (rst) begin // @[tsqr_fsm.scala 261:18]
      dmx0_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 265:31]
    end else begin
      dmx0_mem_enb_reg <= _rd_dmx0_en_T_1 & rd_mem_fst | rd_dmx0_en; // @[tsqr_fsm.scala 272:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx1_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 404:26]
    end else if (rst) begin // @[tsqr_fsm.scala 261:18]
      dmx1_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 266:31]
    end else begin
      dmx1_mem_enb_reg <= mx_cnt[0] & rd_mem_fst | rd_dmx1_en; // @[tsqr_fsm.scala 273:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      rtri_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 405:26]
    end else if (rst) begin // @[tsqr_fsm.scala 261:18]
      rtri_mem_enb_reg <= 1'h0; // @[tsqr_fsm.scala 267:31]
    end else begin
      rtri_mem_enb_reg <= rd_mem_fst | rd_rtri_en; // @[tsqr_fsm.scala 274:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx0_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 406:26]
    end else if (rst) begin // @[tsqr_fsm.scala 329:18]
      dmx0_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 330:31]
    end else begin
      dmx0_mem_ena_reg <= _rd_dmx0_en_T_1 & _yjp_vld_T_16 & tr_cnt < _hh_fi_T_1; // @[tsqr_fsm.scala 334:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx1_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 407:26]
    end else if (rst) begin // @[tsqr_fsm.scala 329:18]
      dmx1_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 331:31]
    end else begin
      dmx1_mem_ena_reg <= mx_cnt[0] & _yjp_vld_T_16 & _dmx0_mem_ena_wire_T_6; // @[tsqr_fsm.scala 335:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      rtri_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 408:26]
    end else if (rst) begin // @[tsqr_fsm.scala 329:18]
      rtri_mem_ena_reg <= 1'h0; // @[tsqr_fsm.scala 332:31]
    end else begin
      rtri_mem_ena_reg <= _yjp_vld_T_16 & _dmx0_mem_ena_wire_T_6; // @[tsqr_fsm.scala 336:31]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx0_mem_addrb_reg <= 5'h0; // @[tsqr_fsm.scala 399:28]
    end else begin
      dmx0_mem_addrb_reg <= dmx0_mem_addrb_wire; // @[tsqr_fsm.scala 415:28]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx1_mem_addrb_reg <= 5'h0; // @[tsqr_fsm.scala 400:28]
    end else begin
      dmx1_mem_addrb_reg <= dmx1_mem_addrb_wire; // @[tsqr_fsm.scala 416:28]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      rtri_mem_addrb_reg <= 5'h0; // @[tsqr_fsm.scala 401:28]
    end else begin
      rtri_mem_addrb_reg <= rtri_mem_addrb_wire; // @[tsqr_fsm.scala 417:28]
    end
    if (rst) begin // @[tsqr_fsm.scala 357:18]
      dmx0_mem_wea_reg <= 128'h0; // @[tsqr_fsm.scala 358:30]
    end else begin
      dmx0_mem_wea_reg <= dmx0_mem_wea; // @[tsqr_fsm.scala 362:30]
    end
    if (rst) begin // @[tsqr_fsm.scala 357:18]
      dmx1_mem_wea_reg <= 128'h0; // @[tsqr_fsm.scala 359:30]
    end else begin
      dmx1_mem_wea_reg <= dmx1_mem_wea; // @[tsqr_fsm.scala 363:30]
    end
    if (rst) begin // @[tsqr_fsm.scala 357:18]
      rtri_mem_wea_reg <= 128'h0; // @[tsqr_fsm.scala 360:30]
    end else begin
      rtri_mem_wea_reg <= rtri_mem_wea; // @[tsqr_fsm.scala 364:30]
    end
    if (rst) begin // @[tsqr_fsm.scala 442:14]
      rtri_mem_wea_update <= 128'hffffffffffffffffffffffffffffffff; // @[tsqr_fsm.scala 446:29]
    end else if (hh_en & tr_cnt == 16'hf9) begin // @[tsqr_fsm.scala 448:55]
      rtri_mem_wea_update <= _rtri_mem_wea_update_T_3; // @[tsqr_fsm.scala 449:29]
    end else begin
      rtri_mem_wea_update <= 128'hffffffffffffffffffffffffffffffff; // @[tsqr_fsm.scala 454:29]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx0_mem_addra_reg <= 5'h0; // @[tsqr_fsm.scala 396:28]
    end else begin
      dmx0_mem_addra_reg <= dmx0_mem_addra_wire; // @[tsqr_fsm.scala 412:28]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      dmx1_mem_addra_reg <= 5'h0; // @[tsqr_fsm.scala 397:28]
    end else begin
      dmx1_mem_addra_reg <= dmx1_mem_addra_wire; // @[tsqr_fsm.scala 413:28]
    end
    if (rst) begin // @[tsqr_fsm.scala 395:14]
      rtri_mem_addra_reg <= 5'h0; // @[tsqr_fsm.scala 398:28]
    end else begin
      rtri_mem_addra_reg <= rtri_mem_addra_wire; // @[tsqr_fsm.scala 414:28]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hh_en = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  nxt_hh_cnt = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  nxt_mx_cnt = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  tr_cy_reg = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  tr_cnt_en = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tr_cnt = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  d1_rdy_REG = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  d1_vld_REG = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  d2_vld_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  vk1_vld_REG = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  d3_rdy_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  d3_vld_REG = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  tk_vld_REG = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  dmx0_mem_enb_reg = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  dmx1_mem_enb_reg = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  rtri_mem_enb_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  dmx0_mem_ena_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  dmx1_mem_ena_reg = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  rtri_mem_ena_reg = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  dmx0_mem_addrb_reg = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  dmx1_mem_addrb_reg = _RAND_21[4:0];
  _RAND_22 = {1{`RANDOM}};
  rtri_mem_addrb_reg = _RAND_22[4:0];
  _RAND_23 = {4{`RANDOM}};
  dmx0_mem_wea_reg = _RAND_23[127:0];
  _RAND_24 = {4{`RANDOM}};
  dmx1_mem_wea_reg = _RAND_24[127:0];
  _RAND_25 = {4{`RANDOM}};
  rtri_mem_wea_reg = _RAND_25[127:0];
  _RAND_26 = {4{`RANDOM}};
  rtri_mem_wea_update = _RAND_26[127:0];
  _RAND_27 = {1{`RANDOM}};
  dmx0_mem_addra_reg = _RAND_27[4:0];
  _RAND_28 = {1{`RANDOM}};
  dmx1_mem_addra_reg = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  rtri_mem_addra_reg = _RAND_29[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module simple_dual(
  input           io_clka,
  input           io_clkb,
  input           io_ena,
  input           io_enb,
  input  [127:0]  io_wea,
  input  [4:0]    io_addra,
  input  [4:0]    io_addrb,
  input  [1023:0] io_dina,
  output [1023:0] io_doutb
);
`ifdef RANDOMIZE_MEM_INIT
  reg [1023:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [1023:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1023:0] ram [0:31]; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_31_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_31_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_31_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_30_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_30_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_30_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_29_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_29_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_29_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_28_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_28_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_28_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_27_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_27_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_27_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_26_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_26_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_26_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_25_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_25_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_25_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_24_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_24_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_24_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_23_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_23_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_23_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_22_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_22_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_22_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_21_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_21_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_21_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_20_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_20_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_20_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_19_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_19_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_19_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_18_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_18_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_18_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_17_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_17_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_17_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_16_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_16_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_16_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_15_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_15_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_15_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_14_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_14_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_14_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_13_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_13_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_13_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_12_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_12_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_12_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_11_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_11_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_11_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_10_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_10_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_10_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_9_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_9_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_9_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_8_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_8_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_8_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_7_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_7_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_7_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_6_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_6_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_6_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_5_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_5_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_5_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_4_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_4_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_4_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_3_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_3_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_3_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_2_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_2_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_2_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_1_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_1_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_1_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_ramtemp_0_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_ramtemp_0_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_ramtemp_0_MPORT_data; // @[hh_core.scala 249:26]
  wire  ram_doutb_MPORT_en; // @[hh_core.scala 249:26]
  wire [4:0] ram_doutb_MPORT_addr; // @[hh_core.scala 249:26]
  wire [1023:0] ram_doutb_MPORT_data; // @[hh_core.scala 249:26]
  wire [1023:0] ram_MPORT_data; // @[hh_core.scala 249:26]
  wire [4:0] ram_MPORT_addr; // @[hh_core.scala 249:26]
  wire  ram_MPORT_mask; // @[hh_core.scala 249:26]
  wire  ram_MPORT_en; // @[hh_core.scala 249:26]
  reg [1023:0] doutb; // @[hh_core.scala 246:28]
  wire [31:0] _dintemp_31_T_9 = {io_wea[127:124],io_wea[127:124],io_wea[127:124],io_wea[127:124],io_wea[127:124],io_wea[
    127:124],io_wea[127:124],io_wea[127:124]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_31_T_10 = io_dina[1023:992] & _dintemp_31_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_31_T_10 = ~_dintemp_31_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_31_T_11 = ram_ramtemp_31_MPORT_data[1023:992] & _ramtemp_31_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_30_T_9 = {io_wea[123:120],io_wea[123:120],io_wea[123:120],io_wea[123:120],io_wea[123:120],io_wea[
    123:120],io_wea[123:120],io_wea[123:120]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_30_T_10 = io_dina[991:960] & _dintemp_30_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_30_T_10 = ~_dintemp_30_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_30_T_11 = ram_ramtemp_30_MPORT_data[991:960] & _ramtemp_30_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_29_T_9 = {io_wea[119:116],io_wea[119:116],io_wea[119:116],io_wea[119:116],io_wea[119:116],io_wea[
    119:116],io_wea[119:116],io_wea[119:116]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_29_T_10 = io_dina[959:928] & _dintemp_29_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_29_T_10 = ~_dintemp_29_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_29_T_11 = ram_ramtemp_29_MPORT_data[959:928] & _ramtemp_29_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_28_T_9 = {io_wea[115:112],io_wea[115:112],io_wea[115:112],io_wea[115:112],io_wea[115:112],io_wea[
    115:112],io_wea[115:112],io_wea[115:112]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_28_T_10 = io_dina[927:896] & _dintemp_28_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_28_T_10 = ~_dintemp_28_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_28_T_11 = ram_ramtemp_28_MPORT_data[927:896] & _ramtemp_28_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_27_T_9 = {io_wea[111:108],io_wea[111:108],io_wea[111:108],io_wea[111:108],io_wea[111:108],io_wea[
    111:108],io_wea[111:108],io_wea[111:108]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_27_T_10 = io_dina[895:864] & _dintemp_27_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_27_T_10 = ~_dintemp_27_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_27_T_11 = ram_ramtemp_27_MPORT_data[895:864] & _ramtemp_27_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_26_T_9 = {io_wea[107:104],io_wea[107:104],io_wea[107:104],io_wea[107:104],io_wea[107:104],io_wea[
    107:104],io_wea[107:104],io_wea[107:104]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_26_T_10 = io_dina[863:832] & _dintemp_26_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_26_T_10 = ~_dintemp_26_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_26_T_11 = ram_ramtemp_26_MPORT_data[863:832] & _ramtemp_26_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_25_T_9 = {io_wea[103:100],io_wea[103:100],io_wea[103:100],io_wea[103:100],io_wea[103:100],io_wea[
    103:100],io_wea[103:100],io_wea[103:100]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_25_T_10 = io_dina[831:800] & _dintemp_25_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_25_T_10 = ~_dintemp_25_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_25_T_11 = ram_ramtemp_25_MPORT_data[831:800] & _ramtemp_25_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_24_T_9 = {io_wea[99:96],io_wea[99:96],io_wea[99:96],io_wea[99:96],io_wea[99:96],io_wea[99:96],
    io_wea[99:96],io_wea[99:96]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_24_T_10 = io_dina[799:768] & _dintemp_24_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_24_T_10 = ~_dintemp_24_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_24_T_11 = ram_ramtemp_24_MPORT_data[799:768] & _ramtemp_24_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_23_T_9 = {io_wea[95:92],io_wea[95:92],io_wea[95:92],io_wea[95:92],io_wea[95:92],io_wea[95:92],
    io_wea[95:92],io_wea[95:92]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_23_T_10 = io_dina[767:736] & _dintemp_23_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_23_T_10 = ~_dintemp_23_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_23_T_11 = ram_ramtemp_23_MPORT_data[767:736] & _ramtemp_23_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_22_T_9 = {io_wea[91:88],io_wea[91:88],io_wea[91:88],io_wea[91:88],io_wea[91:88],io_wea[91:88],
    io_wea[91:88],io_wea[91:88]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_22_T_10 = io_dina[735:704] & _dintemp_22_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_22_T_10 = ~_dintemp_22_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_22_T_11 = ram_ramtemp_22_MPORT_data[735:704] & _ramtemp_22_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_21_T_9 = {io_wea[87:84],io_wea[87:84],io_wea[87:84],io_wea[87:84],io_wea[87:84],io_wea[87:84],
    io_wea[87:84],io_wea[87:84]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_21_T_10 = io_dina[703:672] & _dintemp_21_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_21_T_10 = ~_dintemp_21_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_21_T_11 = ram_ramtemp_21_MPORT_data[703:672] & _ramtemp_21_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_20_T_9 = {io_wea[83:80],io_wea[83:80],io_wea[83:80],io_wea[83:80],io_wea[83:80],io_wea[83:80],
    io_wea[83:80],io_wea[83:80]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_20_T_10 = io_dina[671:640] & _dintemp_20_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_20_T_10 = ~_dintemp_20_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_20_T_11 = ram_ramtemp_20_MPORT_data[671:640] & _ramtemp_20_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_19_T_9 = {io_wea[79:76],io_wea[79:76],io_wea[79:76],io_wea[79:76],io_wea[79:76],io_wea[79:76],
    io_wea[79:76],io_wea[79:76]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_19_T_10 = io_dina[639:608] & _dintemp_19_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_19_T_10 = ~_dintemp_19_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_19_T_11 = ram_ramtemp_19_MPORT_data[639:608] & _ramtemp_19_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_18_T_9 = {io_wea[75:72],io_wea[75:72],io_wea[75:72],io_wea[75:72],io_wea[75:72],io_wea[75:72],
    io_wea[75:72],io_wea[75:72]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_18_T_10 = io_dina[607:576] & _dintemp_18_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_18_T_10 = ~_dintemp_18_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_18_T_11 = ram_ramtemp_18_MPORT_data[607:576] & _ramtemp_18_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_17_T_9 = {io_wea[71:68],io_wea[71:68],io_wea[71:68],io_wea[71:68],io_wea[71:68],io_wea[71:68],
    io_wea[71:68],io_wea[71:68]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_17_T_10 = io_dina[575:544] & _dintemp_17_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_17_T_10 = ~_dintemp_17_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_17_T_11 = ram_ramtemp_17_MPORT_data[575:544] & _ramtemp_17_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_16_T_9 = {io_wea[67:64],io_wea[67:64],io_wea[67:64],io_wea[67:64],io_wea[67:64],io_wea[67:64],
    io_wea[67:64],io_wea[67:64]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_16_T_10 = io_dina[543:512] & _dintemp_16_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_16_T_10 = ~_dintemp_16_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_16_T_11 = ram_ramtemp_16_MPORT_data[543:512] & _ramtemp_16_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_15_T_9 = {io_wea[63:60],io_wea[63:60],io_wea[63:60],io_wea[63:60],io_wea[63:60],io_wea[63:60],
    io_wea[63:60],io_wea[63:60]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_15_T_10 = io_dina[511:480] & _dintemp_15_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_15_T_10 = ~_dintemp_15_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_15_T_11 = ram_ramtemp_15_MPORT_data[511:480] & _ramtemp_15_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_14_T_9 = {io_wea[59:56],io_wea[59:56],io_wea[59:56],io_wea[59:56],io_wea[59:56],io_wea[59:56],
    io_wea[59:56],io_wea[59:56]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_14_T_10 = io_dina[479:448] & _dintemp_14_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_14_T_10 = ~_dintemp_14_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_14_T_11 = ram_ramtemp_14_MPORT_data[479:448] & _ramtemp_14_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_13_T_9 = {io_wea[55:52],io_wea[55:52],io_wea[55:52],io_wea[55:52],io_wea[55:52],io_wea[55:52],
    io_wea[55:52],io_wea[55:52]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_13_T_10 = io_dina[447:416] & _dintemp_13_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_13_T_10 = ~_dintemp_13_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_13_T_11 = ram_ramtemp_13_MPORT_data[447:416] & _ramtemp_13_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_12_T_9 = {io_wea[51:48],io_wea[51:48],io_wea[51:48],io_wea[51:48],io_wea[51:48],io_wea[51:48],
    io_wea[51:48],io_wea[51:48]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_12_T_10 = io_dina[415:384] & _dintemp_12_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_12_T_10 = ~_dintemp_12_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_12_T_11 = ram_ramtemp_12_MPORT_data[415:384] & _ramtemp_12_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_11_T_9 = {io_wea[47:44],io_wea[47:44],io_wea[47:44],io_wea[47:44],io_wea[47:44],io_wea[47:44],
    io_wea[47:44],io_wea[47:44]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_11_T_10 = io_dina[383:352] & _dintemp_11_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_11_T_10 = ~_dintemp_11_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_11_T_11 = ram_ramtemp_11_MPORT_data[383:352] & _ramtemp_11_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_10_T_9 = {io_wea[43:40],io_wea[43:40],io_wea[43:40],io_wea[43:40],io_wea[43:40],io_wea[43:40],
    io_wea[43:40],io_wea[43:40]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_10_T_10 = io_dina[351:320] & _dintemp_10_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_10_T_10 = ~_dintemp_10_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_10_T_11 = ram_ramtemp_10_MPORT_data[351:320] & _ramtemp_10_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_9_T_9 = {io_wea[39:36],io_wea[39:36],io_wea[39:36],io_wea[39:36],io_wea[39:36],io_wea[39:36],
    io_wea[39:36],io_wea[39:36]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_9_T_10 = io_dina[319:288] & _dintemp_9_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_9_T_10 = ~_dintemp_9_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_9_T_11 = ram_ramtemp_9_MPORT_data[319:288] & _ramtemp_9_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_8_T_9 = {io_wea[35:32],io_wea[35:32],io_wea[35:32],io_wea[35:32],io_wea[35:32],io_wea[35:32],
    io_wea[35:32],io_wea[35:32]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_8_T_10 = io_dina[287:256] & _dintemp_8_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_8_T_10 = ~_dintemp_8_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_8_T_11 = ram_ramtemp_8_MPORT_data[287:256] & _ramtemp_8_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_7_T_9 = {io_wea[31:28],io_wea[31:28],io_wea[31:28],io_wea[31:28],io_wea[31:28],io_wea[31:28],
    io_wea[31:28],io_wea[31:28]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_7_T_10 = io_dina[255:224] & _dintemp_7_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_7_T_10 = ~_dintemp_7_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_7_T_11 = ram_ramtemp_7_MPORT_data[255:224] & _ramtemp_7_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_6_T_9 = {io_wea[27:24],io_wea[27:24],io_wea[27:24],io_wea[27:24],io_wea[27:24],io_wea[27:24],
    io_wea[27:24],io_wea[27:24]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_6_T_10 = io_dina[223:192] & _dintemp_6_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_6_T_10 = ~_dintemp_6_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_6_T_11 = ram_ramtemp_6_MPORT_data[223:192] & _ramtemp_6_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_5_T_9 = {io_wea[23:20],io_wea[23:20],io_wea[23:20],io_wea[23:20],io_wea[23:20],io_wea[23:20],
    io_wea[23:20],io_wea[23:20]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_5_T_10 = io_dina[191:160] & _dintemp_5_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_5_T_10 = ~_dintemp_5_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_5_T_11 = ram_ramtemp_5_MPORT_data[191:160] & _ramtemp_5_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_4_T_9 = {io_wea[19:16],io_wea[19:16],io_wea[19:16],io_wea[19:16],io_wea[19:16],io_wea[19:16],
    io_wea[19:16],io_wea[19:16]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_4_T_10 = io_dina[159:128] & _dintemp_4_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_4_T_10 = ~_dintemp_4_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_4_T_11 = ram_ramtemp_4_MPORT_data[159:128] & _ramtemp_4_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_3_T_9 = {io_wea[15:12],io_wea[15:12],io_wea[15:12],io_wea[15:12],io_wea[15:12],io_wea[15:12],
    io_wea[15:12],io_wea[15:12]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_3_T_10 = io_dina[127:96] & _dintemp_3_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_3_T_10 = ~_dintemp_3_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_3_T_11 = ram_ramtemp_3_MPORT_data[127:96] & _ramtemp_3_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_2_T_9 = {io_wea[11:8],io_wea[11:8],io_wea[11:8],io_wea[11:8],io_wea[11:8],io_wea[11:8],io_wea[11:
    8],io_wea[11:8]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_2_T_10 = io_dina[95:64] & _dintemp_2_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_2_T_10 = ~_dintemp_2_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_2_T_11 = ram_ramtemp_2_MPORT_data[95:64] & _ramtemp_2_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_1_T_9 = {io_wea[7:4],io_wea[7:4],io_wea[7:4],io_wea[7:4],io_wea[7:4],io_wea[7:4],io_wea[7:4],
    io_wea[7:4]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_1_T_10 = io_dina[63:32] & _dintemp_1_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_1_T_10 = ~_dintemp_1_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_1_T_11 = ram_ramtemp_1_MPORT_data[63:32] & _ramtemp_1_T_10; // @[hh_core.scala 263:131]
  wire [31:0] _dintemp_0_T_9 = {io_wea[3:0],io_wea[3:0],io_wea[3:0],io_wea[3:0],io_wea[3:0],io_wea[3:0],io_wea[3:0],
    io_wea[3:0]}; // @[Cat.scala 31:58]
  wire [31:0] _dintemp_0_T_10 = io_dina[31:0] & _dintemp_0_T_9; // @[hh_core.scala 259:123]
  wire [31:0] _ramtemp_0_T_10 = ~_dintemp_0_T_9; // @[hh_core.scala 263:133]
  wire [31:0] _ramtemp_0_T_11 = ram_ramtemp_0_MPORT_data[31:0] & _ramtemp_0_T_10; // @[hh_core.scala 263:131]
  wire [31:0] ramtemp_1 = io_ena ? _ramtemp_1_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_0 = io_ena ? _ramtemp_0_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_3 = io_ena ? _ramtemp_3_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_2 = io_ena ? _ramtemp_2_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_5 = io_ena ? _ramtemp_5_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_4 = io_ena ? _ramtemp_4_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_7 = io_ena ? _ramtemp_7_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_6 = io_ena ? _ramtemp_6_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [255:0] lo_lo = {ramtemp_7,ramtemp_6,ramtemp_5,ramtemp_4,ramtemp_3,ramtemp_2,ramtemp_1,ramtemp_0}; // @[hh_core.scala 265:45]
  wire [31:0] ramtemp_9 = io_ena ? _ramtemp_9_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_8 = io_ena ? _ramtemp_8_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_11 = io_ena ? _ramtemp_11_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_10 = io_ena ? _ramtemp_10_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_13 = io_ena ? _ramtemp_13_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_12 = io_ena ? _ramtemp_12_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_15 = io_ena ? _ramtemp_15_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_14 = io_ena ? _ramtemp_14_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [511:0] lo = {ramtemp_15,ramtemp_14,ramtemp_13,ramtemp_12,ramtemp_11,ramtemp_10,ramtemp_9,ramtemp_8,lo_lo}; // @[hh_core.scala 265:45]
  wire [31:0] ramtemp_17 = io_ena ? _ramtemp_17_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_16 = io_ena ? _ramtemp_16_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_19 = io_ena ? _ramtemp_19_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_18 = io_ena ? _ramtemp_18_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_21 = io_ena ? _ramtemp_21_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_20 = io_ena ? _ramtemp_20_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_23 = io_ena ? _ramtemp_23_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_22 = io_ena ? _ramtemp_22_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [255:0] hi_lo = {ramtemp_23,ramtemp_22,ramtemp_21,ramtemp_20,ramtemp_19,ramtemp_18,ramtemp_17,ramtemp_16}; // @[hh_core.scala 265:45]
  wire [31:0] ramtemp_25 = io_ena ? _ramtemp_25_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_24 = io_ena ? _ramtemp_24_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_27 = io_ena ? _ramtemp_27_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_26 = io_ena ? _ramtemp_26_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_29 = io_ena ? _ramtemp_29_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_28 = io_ena ? _ramtemp_28_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_31 = io_ena ? _ramtemp_31_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [31:0] ramtemp_30 = io_ena ? _ramtemp_30_T_11 : 32'h0; // @[hh_core.scala 255:25 263:48 269:28]
  wire [1023:0] _T = {ramtemp_31,ramtemp_30,ramtemp_29,ramtemp_28,ramtemp_27,ramtemp_26,ramtemp_25,ramtemp_24,hi_lo,lo}; // @[hh_core.scala 265:45]
  wire [31:0] dintemp_1 = io_ena ? _dintemp_1_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_0 = io_ena ? _dintemp_0_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_3 = io_ena ? _dintemp_3_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_2 = io_ena ? _dintemp_2_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_5 = io_ena ? _dintemp_5_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_4 = io_ena ? _dintemp_4_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_7 = io_ena ? _dintemp_7_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_6 = io_ena ? _dintemp_6_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [255:0] lo_lo_1 = {dintemp_7,dintemp_6,dintemp_5,dintemp_4,dintemp_3,dintemp_2,dintemp_1,dintemp_0}; // @[hh_core.scala 265:62]
  wire [31:0] dintemp_9 = io_ena ? _dintemp_9_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_8 = io_ena ? _dintemp_8_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_11 = io_ena ? _dintemp_11_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_10 = io_ena ? _dintemp_10_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_13 = io_ena ? _dintemp_13_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_12 = io_ena ? _dintemp_12_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_15 = io_ena ? _dintemp_15_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_14 = io_ena ? _dintemp_14_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [511:0] lo_1 = {dintemp_15,dintemp_14,dintemp_13,dintemp_12,dintemp_11,dintemp_10,dintemp_9,dintemp_8,lo_lo_1}; // @[hh_core.scala 265:62]
  wire [31:0] dintemp_17 = io_ena ? _dintemp_17_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_16 = io_ena ? _dintemp_16_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_19 = io_ena ? _dintemp_19_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_18 = io_ena ? _dintemp_18_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_21 = io_ena ? _dintemp_21_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_20 = io_ena ? _dintemp_20_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_23 = io_ena ? _dintemp_23_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_22 = io_ena ? _dintemp_22_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [255:0] hi_lo_1 = {dintemp_23,dintemp_22,dintemp_21,dintemp_20,dintemp_19,dintemp_18,dintemp_17,dintemp_16}; // @[hh_core.scala 265:62]
  wire [31:0] dintemp_25 = io_ena ? _dintemp_25_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_24 = io_ena ? _dintemp_24_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_27 = io_ena ? _dintemp_27_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_26 = io_ena ? _dintemp_26_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_29 = io_ena ? _dintemp_29_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_28 = io_ena ? _dintemp_28_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_31 = io_ena ? _dintemp_31_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [31:0] dintemp_30 = io_ena ? _dintemp_30_T_10 : 32'h0; // @[hh_core.scala 255:25 259:48 268:28]
  wire [1023:0] _T_1 = {dintemp_31,dintemp_30,dintemp_29,dintemp_28,dintemp_27,dintemp_26,dintemp_25,dintemp_24,hi_lo_1,
    lo_1}; // @[hh_core.scala 265:62]
  assign ram_ramtemp_31_MPORT_en = io_ena;
  assign ram_ramtemp_31_MPORT_addr = io_addra;
  assign ram_ramtemp_31_MPORT_data = ram[ram_ramtemp_31_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_30_MPORT_en = io_ena;
  assign ram_ramtemp_30_MPORT_addr = io_addra;
  assign ram_ramtemp_30_MPORT_data = ram[ram_ramtemp_30_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_29_MPORT_en = io_ena;
  assign ram_ramtemp_29_MPORT_addr = io_addra;
  assign ram_ramtemp_29_MPORT_data = ram[ram_ramtemp_29_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_28_MPORT_en = io_ena;
  assign ram_ramtemp_28_MPORT_addr = io_addra;
  assign ram_ramtemp_28_MPORT_data = ram[ram_ramtemp_28_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_27_MPORT_en = io_ena;
  assign ram_ramtemp_27_MPORT_addr = io_addra;
  assign ram_ramtemp_27_MPORT_data = ram[ram_ramtemp_27_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_26_MPORT_en = io_ena;
  assign ram_ramtemp_26_MPORT_addr = io_addra;
  assign ram_ramtemp_26_MPORT_data = ram[ram_ramtemp_26_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_25_MPORT_en = io_ena;
  assign ram_ramtemp_25_MPORT_addr = io_addra;
  assign ram_ramtemp_25_MPORT_data = ram[ram_ramtemp_25_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_24_MPORT_en = io_ena;
  assign ram_ramtemp_24_MPORT_addr = io_addra;
  assign ram_ramtemp_24_MPORT_data = ram[ram_ramtemp_24_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_23_MPORT_en = io_ena;
  assign ram_ramtemp_23_MPORT_addr = io_addra;
  assign ram_ramtemp_23_MPORT_data = ram[ram_ramtemp_23_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_22_MPORT_en = io_ena;
  assign ram_ramtemp_22_MPORT_addr = io_addra;
  assign ram_ramtemp_22_MPORT_data = ram[ram_ramtemp_22_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_21_MPORT_en = io_ena;
  assign ram_ramtemp_21_MPORT_addr = io_addra;
  assign ram_ramtemp_21_MPORT_data = ram[ram_ramtemp_21_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_20_MPORT_en = io_ena;
  assign ram_ramtemp_20_MPORT_addr = io_addra;
  assign ram_ramtemp_20_MPORT_data = ram[ram_ramtemp_20_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_19_MPORT_en = io_ena;
  assign ram_ramtemp_19_MPORT_addr = io_addra;
  assign ram_ramtemp_19_MPORT_data = ram[ram_ramtemp_19_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_18_MPORT_en = io_ena;
  assign ram_ramtemp_18_MPORT_addr = io_addra;
  assign ram_ramtemp_18_MPORT_data = ram[ram_ramtemp_18_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_17_MPORT_en = io_ena;
  assign ram_ramtemp_17_MPORT_addr = io_addra;
  assign ram_ramtemp_17_MPORT_data = ram[ram_ramtemp_17_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_16_MPORT_en = io_ena;
  assign ram_ramtemp_16_MPORT_addr = io_addra;
  assign ram_ramtemp_16_MPORT_data = ram[ram_ramtemp_16_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_15_MPORT_en = io_ena;
  assign ram_ramtemp_15_MPORT_addr = io_addra;
  assign ram_ramtemp_15_MPORT_data = ram[ram_ramtemp_15_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_14_MPORT_en = io_ena;
  assign ram_ramtemp_14_MPORT_addr = io_addra;
  assign ram_ramtemp_14_MPORT_data = ram[ram_ramtemp_14_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_13_MPORT_en = io_ena;
  assign ram_ramtemp_13_MPORT_addr = io_addra;
  assign ram_ramtemp_13_MPORT_data = ram[ram_ramtemp_13_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_12_MPORT_en = io_ena;
  assign ram_ramtemp_12_MPORT_addr = io_addra;
  assign ram_ramtemp_12_MPORT_data = ram[ram_ramtemp_12_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_11_MPORT_en = io_ena;
  assign ram_ramtemp_11_MPORT_addr = io_addra;
  assign ram_ramtemp_11_MPORT_data = ram[ram_ramtemp_11_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_10_MPORT_en = io_ena;
  assign ram_ramtemp_10_MPORT_addr = io_addra;
  assign ram_ramtemp_10_MPORT_data = ram[ram_ramtemp_10_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_9_MPORT_en = io_ena;
  assign ram_ramtemp_9_MPORT_addr = io_addra;
  assign ram_ramtemp_9_MPORT_data = ram[ram_ramtemp_9_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_8_MPORT_en = io_ena;
  assign ram_ramtemp_8_MPORT_addr = io_addra;
  assign ram_ramtemp_8_MPORT_data = ram[ram_ramtemp_8_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_7_MPORT_en = io_ena;
  assign ram_ramtemp_7_MPORT_addr = io_addra;
  assign ram_ramtemp_7_MPORT_data = ram[ram_ramtemp_7_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_6_MPORT_en = io_ena;
  assign ram_ramtemp_6_MPORT_addr = io_addra;
  assign ram_ramtemp_6_MPORT_data = ram[ram_ramtemp_6_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_5_MPORT_en = io_ena;
  assign ram_ramtemp_5_MPORT_addr = io_addra;
  assign ram_ramtemp_5_MPORT_data = ram[ram_ramtemp_5_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_4_MPORT_en = io_ena;
  assign ram_ramtemp_4_MPORT_addr = io_addra;
  assign ram_ramtemp_4_MPORT_data = ram[ram_ramtemp_4_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_3_MPORT_en = io_ena;
  assign ram_ramtemp_3_MPORT_addr = io_addra;
  assign ram_ramtemp_3_MPORT_data = ram[ram_ramtemp_3_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_2_MPORT_en = io_ena;
  assign ram_ramtemp_2_MPORT_addr = io_addra;
  assign ram_ramtemp_2_MPORT_data = ram[ram_ramtemp_2_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_1_MPORT_en = io_ena;
  assign ram_ramtemp_1_MPORT_addr = io_addra;
  assign ram_ramtemp_1_MPORT_data = ram[ram_ramtemp_1_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_ramtemp_0_MPORT_en = io_ena;
  assign ram_ramtemp_0_MPORT_addr = io_addra;
  assign ram_ramtemp_0_MPORT_data = ram[ram_ramtemp_0_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_doutb_MPORT_en = io_enb;
  assign ram_doutb_MPORT_addr = io_addrb;
  assign ram_doutb_MPORT_data = ram[ram_doutb_MPORT_addr]; // @[hh_core.scala 249:26]
  assign ram_MPORT_data = _T + _T_1;
  assign ram_MPORT_addr = io_addra;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_ena;
  assign io_doutb = doutb; // @[hh_core.scala 247:22]
  always @(posedge io_clka) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[hh_core.scala 249:26]
    end
    if (io_enb) begin // @[hh_core.scala 273:29]
      doutb <= ram_doutb_MPORT_data; // @[hh_core.scala 274:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {32{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[1023:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {32{`RANDOM}};
  doutb = _RAND_1[1023:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module multiplier(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [47:0] io_out_s
);
  assign io_out_s = io_in_a * io_in_b; // @[BinaryDesigns.scala 81:23]
endmodule
module full_subber(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a - io_in_b; // @[BinaryDesigns.scala 69:23]
  wire [9:0] _result_T_2 = _result_T - 9'h0; // @[BinaryDesigns.scala 69:34]
  wire [8:0] result = _result_T_2[8:0]; // @[BinaryDesigns.scala 68:22 69:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 70:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 71:23]
endmodule
module twoscomplement(
  input  [7:0] io_in,
  output [7:0] io_out
);
  wire [7:0] _x_T = ~io_in; // @[BinaryDesigns.scala 25:16]
  assign io_out = 8'h1 + _x_T; // @[BinaryDesigns.scala 25:14]
endmodule
module full_adder(
  input  [7:0] io_in_a,
  input  [7:0] io_in_b,
  output [7:0] io_out_s,
  output       io_out_c
);
  wire [8:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [9:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [8:0] result = _result_T_1[8:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[7:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[8]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_multiplier_10ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] multiplier_io_in_a; // @[FloatingPointDesigns.scala 1723:28]
  wire [23:0] multiplier_io_in_b; // @[FloatingPointDesigns.scala 1723:28]
  wire [47:0] multiplier_io_out_s; // @[FloatingPointDesigns.scala 1723:28]
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1730:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1730:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1730:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1730:24]
  wire [7:0] complementN_io_in; // @[FloatingPointDesigns.scala 1739:29]
  wire [7:0] complementN_io_out; // @[FloatingPointDesigns.scala 1739:29]
  wire [7:0] adderN_io_in_a; // @[FloatingPointDesigns.scala 1756:24]
  wire [7:0] adderN_io_in_b; // @[FloatingPointDesigns.scala 1756:24]
  wire [7:0] adderN_io_out_s; // @[FloatingPointDesigns.scala 1756:24]
  wire  adderN_io_out_c; // @[FloatingPointDesigns.scala 1756:24]
  wire  s_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1689:20]
  wire  s_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1690:20]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1694:64]
  wire [8:0] _GEN_63 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1694:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1696:45 1697:14 1699:14]
  wire [8:0] _GEN_1 = _GEN_63 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1694:71 1695:14]
  wire [8:0] _GEN_64 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1701:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1703:45 1704:14 1706:14]
  wire [8:0] _GEN_3 = _GEN_64 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1701:71 1702:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1711:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1712:23]
  wire [23:0] new_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1716:24]
  wire [23:0] new_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1717:24]
  reg  s_reg_0_0; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_0_1; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_1_0; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_1_1; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_2_0; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_2_1; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_3_0; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_3_1; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_4_0; // @[FloatingPointDesigns.scala 1719:24]
  reg  s_reg_4_1; // @[FloatingPointDesigns.scala 1719:24]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_3_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_3_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_4_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_4_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_5_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_5_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_6_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_6_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_7_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_7_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_8_0; // @[FloatingPointDesigns.scala 1720:26]
  reg [7:0] exp_reg_8_1; // @[FloatingPointDesigns.scala 1720:26]
  reg [23:0] new_frac_reg_0_0; // @[FloatingPointDesigns.scala 1721:31]
  reg [23:0] new_frac_reg_0_1; // @[FloatingPointDesigns.scala 1721:31]
  reg [23:0] new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1721:31]
  reg [23:0] new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1721:31]
  reg [47:0] multipplier_out_s_reg_0; // @[FloatingPointDesigns.scala 1727:40]
  reg [47:0] multipplier_out_s_reg_1; // @[FloatingPointDesigns.scala 1727:40]
  reg [47:0] multipplier_out_s_reg_2; // @[FloatingPointDesigns.scala 1727:40]
  reg [47:0] multipplier_out_s_reg_3; // @[FloatingPointDesigns.scala 1727:40]
  reg [47:0] multipplier_out_s_reg_4; // @[FloatingPointDesigns.scala 1727:40]
  reg [47:0] multipplier_out_s_reg_5; // @[FloatingPointDesigns.scala 1727:40]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1735:35]
  reg [7:0] complementN_out_reg_0; // @[FloatingPointDesigns.scala 1742:38]
  reg [7:0] complementN_out_reg_1; // @[FloatingPointDesigns.scala 1742:38]
  reg [7:0] complementN_out_reg_2; // @[FloatingPointDesigns.scala 1742:38]
  wire  new_s = s_reg_4_0 ^ s_reg_4_1; // @[FloatingPointDesigns.scala 1745:26]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1747:28]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1747:28]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1747:28]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1747:28]
  wire  is_exp1_neg_wire = exp_reg_5_1 < 8'h7f; // @[FloatingPointDesigns.scala 1750:40]
  reg  is_exp1_neg_reg_0; // @[FloatingPointDesigns.scala 1752:34]
  reg  is_exp1_neg_reg_1; // @[FloatingPointDesigns.scala 1752:34]
  wire [7:0] _adderN_io_in_a_T_1 = exp_reg_6_0 + 8'h1; // @[FloatingPointDesigns.scala 1760:39]
  reg [7:0] adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1767:35]
  reg  adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1768:35]
  reg [7:0] new_exp_reg_0; // @[FloatingPointDesigns.scala 1770:30]
  reg [22:0] new_mant_reg_0; // @[FloatingPointDesigns.scala 1771:31]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1773:28]
  wire  _new_exp_reg_0_T_1 = ~adderN_out_c_reg_0; // @[FloatingPointDesigns.scala 1777:55]
  wire [7:0] _new_exp_reg_0_T_2 = ~adderN_out_c_reg_0 ? 8'h1 : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1777:54]
  wire  _new_exp_reg_0_T_5 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe; // @[FloatingPointDesigns.scala 1777:142]
  wire [7:0] _new_exp_reg_0_T_6 = adderN_out_c_reg_0 | adderN_out_s_reg_0 > 8'hfe ? 8'hfe : adderN_out_s_reg_0; // @[FloatingPointDesigns.scala 1777:114]
  wire [7:0] _new_exp_reg_0_T_7 = is_exp1_neg_reg_1 ? _new_exp_reg_0_T_2 : _new_exp_reg_0_T_6; // @[FloatingPointDesigns.scala 1777:30]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_3,new_exp_reg_0,new_mant_reg_0}; // @[FloatingPointDesigns.scala 1819:53]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1693:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1693:19]
  wire [47:0] _GEN_17 = multiplier_io_out_s; // @[FloatingPointDesigns.scala 1775:19 1787:32 1727:40]
  wire [7:0] _GEN_18 = subber_io_out_s; // @[FloatingPointDesigns.scala 1775:19 1788:27 1735:35]
  wire [7:0] _GEN_20 = complementN_io_out; // @[FloatingPointDesigns.scala 1775:19 1790:30 1742:38]
  wire [7:0] _GEN_23 = adderN_io_out_s; // @[FloatingPointDesigns.scala 1775:19 1793:27 1767:35]
  wire  _GEN_24 = adderN_io_out_c; // @[FloatingPointDesigns.scala 1775:19 1794:27 1768:35]
  multiplier multiplier ( // @[FloatingPointDesigns.scala 1723:28]
    .io_in_a(multiplier_io_in_a),
    .io_in_b(multiplier_io_in_b),
    .io_out_s(multiplier_io_out_s)
  );
  full_subber subber ( // @[FloatingPointDesigns.scala 1730:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  twoscomplement complementN ( // @[FloatingPointDesigns.scala 1739:29]
    .io_in(complementN_io_in),
    .io_out(complementN_io_out)
  );
  full_adder adderN ( // @[FloatingPointDesigns.scala 1756:24]
    .io_in_a(adderN_io_in_a),
    .io_in_b(adderN_io_in_b),
    .io_out_s(adderN_io_out_s),
    .io_out_c(adderN_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1822:14]
  assign multiplier_io_in_a = new_frac_reg_1_0; // @[FloatingPointDesigns.scala 1724:24]
  assign multiplier_io_in_b = new_frac_reg_1_1; // @[FloatingPointDesigns.scala 1725:24]
  assign subber_io_in_a = 8'h7f; // @[FloatingPointDesigns.scala 1731:20]
  assign subber_io_in_b = exp_reg_2_1; // @[FloatingPointDesigns.scala 1732:20]
  assign complementN_io_in = subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1740:23]
  assign adderN_io_in_a = multipplier_out_s_reg_4[47] ? _adderN_io_in_a_T_1 : exp_reg_6_0; // @[FloatingPointDesigns.scala 1759:70 1760:22 1763:22]
  assign adderN_io_in_b = complementN_out_reg_2; // @[FloatingPointDesigns.scala 1759:70 1761:22 1764:22]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_0_0 <= s_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_0_1 <= s_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_1_0 <= s_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_1_1 <= s_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_2_0 <= s_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_2_1 <= s_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_3_0 <= s_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_3_1 <= s_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_4_0 <= s_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1719:24]
      s_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1719:24]
    end else begin
      s_reg_4_1 <= s_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_0_0 <= exp_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_0_1 <= exp_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_1_0 <= exp_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_1_1 <= exp_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_2_0 <= exp_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_2_1 <= exp_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_3_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_3_0 <= exp_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_3_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_3_1 <= exp_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_4_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_4_0 <= exp_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_4_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_4_1 <= exp_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_5_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_5_0 <= exp_reg_4_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_5_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_5_1 <= exp_reg_4_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_6_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_6_0 <= exp_reg_5_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_6_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_6_1 <= exp_reg_5_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_7_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_7_0 <= exp_reg_6_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_7_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_7_1 <= exp_reg_6_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_8_0 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_8_0 <= exp_reg_7_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1720:26]
      exp_reg_8_1 <= 8'h0; // @[FloatingPointDesigns.scala 1720:26]
    end else begin
      exp_reg_8_1 <= exp_reg_7_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1721:31]
      new_frac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1721:31]
    end else begin
      new_frac_reg_0_0 <= new_frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1721:31]
      new_frac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1721:31]
    end else begin
      new_frac_reg_0_1 <= new_frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1721:31]
      new_frac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1721:31]
    end else begin
      new_frac_reg_1_0 <= new_frac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1721:31]
      new_frac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1721:31]
    end else begin
      new_frac_reg_1_1 <= new_frac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_0 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_0 <= _GEN_17;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_1 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_1 <= multipplier_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_2 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_2 <= multipplier_out_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_3 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_3 <= multipplier_out_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_4 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_4 <= multipplier_out_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1727:40]
      multipplier_out_s_reg_5 <= 48'h0; // @[FloatingPointDesigns.scala 1727:40]
    end else begin
      multipplier_out_s_reg_5 <= multipplier_out_s_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1735:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1735:35]
    end else begin
      subber_out_s_reg_0 <= _GEN_18;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1742:38]
      complementN_out_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1742:38]
    end else begin
      complementN_out_reg_0 <= _GEN_20;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1742:38]
      complementN_out_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1742:38]
    end else begin
      complementN_out_reg_1 <= complementN_out_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1742:38]
      complementN_out_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1742:38]
    end else begin
      complementN_out_reg_2 <= complementN_out_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1747:28]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1747:28]
    end else begin
      new_s_reg_0 <= new_s;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1747:28]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1747:28]
    end else begin
      new_s_reg_1 <= new_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1747:28]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1747:28]
    end else begin
      new_s_reg_2 <= new_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1747:28]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1747:28]
    end else begin
      new_s_reg_3 <= new_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1752:34]
      is_exp1_neg_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1752:34]
    end else begin
      is_exp1_neg_reg_0 <= is_exp1_neg_wire;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1752:34]
      is_exp1_neg_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1752:34]
    end else begin
      is_exp1_neg_reg_1 <= is_exp1_neg_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1767:35]
      adderN_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1767:35]
    end else begin
      adderN_out_s_reg_0 <= _GEN_23;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1768:35]
      adderN_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1768:35]
    end else begin
      adderN_out_c_reg_0 <= _GEN_24;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1770:30]
      new_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1770:30]
    end else if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1776:72]
      new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1777:24]
    end else begin
      new_exp_reg_0 <= _new_exp_reg_0_T_7; // @[FloatingPointDesigns.scala 1780:24]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1771:31]
      new_mant_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1771:31]
    end else if (multipplier_out_s_reg_5[47]) begin // @[FloatingPointDesigns.scala 1776:72]
      if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1778:31]
        if (_new_exp_reg_0_T_1) begin // @[FloatingPointDesigns.scala 1778:55]
          new_mant_reg_0 <= 23'h0;
        end else begin
          new_mant_reg_0 <= multipplier_out_s_reg_5[46:24];
        end
      end else if (_new_exp_reg_0_T_5) begin // @[FloatingPointDesigns.scala 1778:160]
        new_mant_reg_0 <= 23'h7fffff;
      end else begin
        new_mant_reg_0 <= multipplier_out_s_reg_5[46:24];
      end
    end else if (is_exp1_neg_reg_1) begin // @[FloatingPointDesigns.scala 1781:31]
      if (_new_exp_reg_0_T_1) begin // @[FloatingPointDesigns.scala 1781:55]
        new_mant_reg_0 <= 23'h0;
      end else begin
        new_mant_reg_0 <= multipplier_out_s_reg_5[45:23];
      end
    end else if (_new_exp_reg_0_T_5) begin // @[FloatingPointDesigns.scala 1781:156]
      new_mant_reg_0 <= 23'h7fffff;
    end else begin
      new_mant_reg_0 <= multipplier_out_s_reg_5[45:23];
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1773:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1773:28]
    end else if (exp_reg_8_0 == 8'h0 | exp_reg_8_1 == 8'h0) begin // @[FloatingPointDesigns.scala 1816:60]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1817:19]
    end else begin
      reg_out_s <= _reg_out_s_T_1; // @[FloatingPointDesigns.scala 1819:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  s_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  s_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  s_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  s_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  s_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  s_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  s_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  s_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  s_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  exp_reg_3_0 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  exp_reg_3_1 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  exp_reg_4_0 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  exp_reg_4_1 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  exp_reg_5_0 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  exp_reg_5_1 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_6_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_6_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_7_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_7_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_8_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_8_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  new_frac_reg_0_0 = _RAND_28[23:0];
  _RAND_29 = {1{`RANDOM}};
  new_frac_reg_0_1 = _RAND_29[23:0];
  _RAND_30 = {1{`RANDOM}};
  new_frac_reg_1_0 = _RAND_30[23:0];
  _RAND_31 = {1{`RANDOM}};
  new_frac_reg_1_1 = _RAND_31[23:0];
  _RAND_32 = {2{`RANDOM}};
  multipplier_out_s_reg_0 = _RAND_32[47:0];
  _RAND_33 = {2{`RANDOM}};
  multipplier_out_s_reg_1 = _RAND_33[47:0];
  _RAND_34 = {2{`RANDOM}};
  multipplier_out_s_reg_2 = _RAND_34[47:0];
  _RAND_35 = {2{`RANDOM}};
  multipplier_out_s_reg_3 = _RAND_35[47:0];
  _RAND_36 = {2{`RANDOM}};
  multipplier_out_s_reg_4 = _RAND_36[47:0];
  _RAND_37 = {2{`RANDOM}};
  multipplier_out_s_reg_5 = _RAND_37[47:0];
  _RAND_38 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  complementN_out_reg_0 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  complementN_out_reg_1 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  complementN_out_reg_2 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  is_exp1_neg_reg_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  is_exp1_neg_reg_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  adderN_out_s_reg_0 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  adderN_out_c_reg_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  new_exp_reg_0 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  new_mant_reg_0 = _RAND_51[22:0];
  _RAND_52 = {1{`RANDOM}};
  reg_out_s = _RAND_52[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module full_adder_64(
  input  [23:0] io_in_a,
  input  [23:0] io_in_b,
  output [23:0] io_out_s,
  output        io_out_c
);
  wire [24:0] _result_T = io_in_a + io_in_b; // @[BinaryDesigns.scala 55:23]
  wire [25:0] _result_T_1 = {{1'd0}, _result_T}; // @[BinaryDesigns.scala 55:34]
  wire [24:0] result = _result_T_1[24:0]; // @[BinaryDesigns.scala 54:22 55:12]
  assign io_out_s = result[23:0]; // @[BinaryDesigns.scala 56:23]
  assign io_out_c = result[24]; // @[BinaryDesigns.scala 57:23]
endmodule
module FP_adder_13ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] subber_io_in_a; // @[FloatingPointDesigns.scala 1456:24]
  wire [7:0] subber_io_in_b; // @[FloatingPointDesigns.scala 1456:24]
  wire [7:0] subber_io_out_s; // @[FloatingPointDesigns.scala 1456:24]
  wire  subber_io_out_c; // @[FloatingPointDesigns.scala 1456:24]
  wire [23:0] adder_io_in_a; // @[FloatingPointDesigns.scala 1462:23]
  wire [23:0] adder_io_in_b; // @[FloatingPointDesigns.scala 1462:23]
  wire [23:0] adder_io_out_s; // @[FloatingPointDesigns.scala 1462:23]
  wire  adder_io_out_c; // @[FloatingPointDesigns.scala 1462:23]
  wire [7:0] subber2_io_in_a; // @[FloatingPointDesigns.scala 1523:25]
  wire [7:0] subber2_io_in_b; // @[FloatingPointDesigns.scala 1523:25]
  wire [7:0] subber2_io_out_s; // @[FloatingPointDesigns.scala 1523:25]
  wire  subber2_io_out_c; // @[FloatingPointDesigns.scala 1523:25]
  wire  sign_0 = io_in_a[31]; // @[FloatingPointDesigns.scala 1385:23]
  wire  sign_1 = io_in_b[31]; // @[FloatingPointDesigns.scala 1386:23]
  wire [8:0] _T_2 = 9'h100 - 9'h2; // @[FloatingPointDesigns.scala 1389:64]
  wire [8:0] _GEN_167 = {{1'd0}, io_in_a[30:23]}; // @[FloatingPointDesigns.scala 1389:36]
  wire [7:0] _GEN_0 = io_in_a[30:23] < 8'h1 ? 8'h1 : io_in_a[30:23]; // @[FloatingPointDesigns.scala 1391:46 1392:14 1394:14]
  wire [8:0] _GEN_1 = _GEN_167 > _T_2 ? _T_2 : {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1389:71 1390:14]
  wire [8:0] _GEN_168 = {{1'd0}, io_in_b[30:23]}; // @[FloatingPointDesigns.scala 1396:36]
  wire [7:0] _GEN_2 = io_in_b[30:23] < 8'h1 ? 8'h1 : io_in_b[30:23]; // @[FloatingPointDesigns.scala 1398:45 1399:14 1401:14]
  wire [8:0] _GEN_3 = _GEN_168 > _T_2 ? _T_2 : {{1'd0}, _GEN_2}; // @[FloatingPointDesigns.scala 1396:71 1397:14]
  wire [22:0] frac_0 = io_in_a[22:0]; // @[FloatingPointDesigns.scala 1406:23]
  wire [22:0] frac_1 = io_in_b[22:0]; // @[FloatingPointDesigns.scala 1407:23]
  wire [23:0] whole_frac_0 = {1'h1,frac_0}; // @[FloatingPointDesigns.scala 1411:26]
  wire [23:0] whole_frac_1 = {1'h1,frac_1}; // @[FloatingPointDesigns.scala 1412:26]
  reg  sign_reg_0_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_0_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_1_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_1_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_2_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_2_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_3_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_3_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_4_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_4_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_5_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_5_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_6_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_6_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_7_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_7_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_8_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_8_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_9_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_9_1; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_10_0; // @[FloatingPointDesigns.scala 1414:28]
  reg  sign_reg_10_1; // @[FloatingPointDesigns.scala 1414:28]
  reg [7:0] exp_reg_0_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_0_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_1_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_1_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_2_0; // @[FloatingPointDesigns.scala 1415:28]
  reg [7:0] exp_reg_2_1; // @[FloatingPointDesigns.scala 1415:28]
  reg [22:0] frac_reg_0_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_0_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_1_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_1_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_2_0; // @[FloatingPointDesigns.scala 1416:28]
  reg [22:0] frac_reg_2_1; // @[FloatingPointDesigns.scala 1416:28]
  reg [23:0] wfrac_reg_0_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_0_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_1_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_1_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1417:28]
  reg [23:0] wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1417:28]
  reg [7:0] subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1419:35]
  reg [7:0] subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1419:35]
  reg  subber_out_c_reg_0; // @[FloatingPointDesigns.scala 1420:35]
  reg  subber_out_c_reg_1; // @[FloatingPointDesigns.scala 1420:35]
  reg [23:0] wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1422:39]
  reg [23:0] wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1422:39]
  reg  ref_s_reg_0; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_1; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_2; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_3; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_4; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_5; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_6; // @[FloatingPointDesigns.scala 1424:31]
  reg  ref_s_reg_7; // @[FloatingPointDesigns.scala 1424:31]
  reg [22:0] ref_frac_reg_0; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_1; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_2; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_3; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_4; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_5; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_6; // @[FloatingPointDesigns.scala 1425:31]
  reg [22:0] ref_frac_reg_7; // @[FloatingPointDesigns.scala 1425:31]
  reg [7:0] ref_exp_reg_0; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_1; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_2; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_3; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_4; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_5; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_6; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] ref_exp_reg_7; // @[FloatingPointDesigns.scala 1426:31]
  reg [7:0] sub_exp_reg_0; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_1; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_2; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_3; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_4; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_5; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_6; // @[FloatingPointDesigns.scala 1427:31]
  reg [7:0] sub_exp_reg_7; // @[FloatingPointDesigns.scala 1427:31]
  reg [23:0] adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1429:37]
  reg [23:0] adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1429:37]
  reg [23:0] adder_io_out_s_reg_2; // @[FloatingPointDesigns.scala 1429:37]
  reg  adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1430:37]
  reg  new_s_reg_0; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_1; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_2; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_3; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_4; // @[FloatingPointDesigns.scala 1432:35]
  reg  new_s_reg_5; // @[FloatingPointDesigns.scala 1432:35]
  reg [22:0] new_out_frac_reg_0; // @[FloatingPointDesigns.scala 1433:35]
  reg [7:0] new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1434:35]
  reg  E_reg_0; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_1; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_2; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_3; // @[FloatingPointDesigns.scala 1435:24]
  reg  E_reg_4; // @[FloatingPointDesigns.scala 1435:24]
  reg  D_reg_0; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_1; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_2; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_3; // @[FloatingPointDesigns.scala 1436:24]
  reg  D_reg_4; // @[FloatingPointDesigns.scala 1436:24]
  reg [23:0] adder_result_reg_0; // @[FloatingPointDesigns.scala 1438:35]
  reg [23:0] adder_result_reg_1; // @[FloatingPointDesigns.scala 1438:35]
  reg [23:0] adder_result_reg_2; // @[FloatingPointDesigns.scala 1438:35]
  reg [5:0] leadingOne_reg_0; // @[FloatingPointDesigns.scala 1440:33]
  reg [5:0] leadingOne_reg_1; // @[FloatingPointDesigns.scala 1440:33]
  reg [31:0] io_in_a_reg_0; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_1; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_2; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_3; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_4; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_5; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_6; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_7; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_8; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_9; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_a_reg_10; // @[FloatingPointDesigns.scala 1442:30]
  reg [31:0] io_in_b_reg_0; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_1; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_2; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_3; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_4; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_5; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_6; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_7; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_8; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_9; // @[FloatingPointDesigns.scala 1443:30]
  reg [31:0] io_in_b_reg_10; // @[FloatingPointDesigns.scala 1443:30]
  reg [7:0] subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1445:36]
  reg  subber2_out_c_reg_0; // @[FloatingPointDesigns.scala 1446:36]
  reg [7:0] cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1467:40]
  wire [7:0] _cmpl_subber_out_s_reg_0_T = ~subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1469:41]
  wire [7:0] _cmpl_subber_out_s_reg_0_T_2 = 8'h1 + _cmpl_subber_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1469:39]
  wire [23:0] _wire_temp_add_in_0_T = wfrac_reg_2_0 >> cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1477:46]
  wire [23:0] _wire_temp_add_in_1_T = wfrac_reg_2_1 >> subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1485:46]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1488:44]
  reg [23:0] cmpl_wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1488:44]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T = ~wire_temp_add_in_reg_0_0; // @[FloatingPointDesigns.scala 1490:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_0_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_0_T; // @[FloatingPointDesigns.scala 1490:46]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T = ~wire_temp_add_in_reg_0_1; // @[FloatingPointDesigns.scala 1491:48]
  wire [23:0] _cmpl_wire_temp_add_in_reg_0_1_T_2 = 24'h1 + _cmpl_wire_temp_add_in_reg_0_1_T; // @[FloatingPointDesigns.scala 1491:46]
  wire [1:0] _adder_io_in_a_T = {sign_reg_4_1,sign_reg_4_0}; // @[FloatingPointDesigns.scala 1494:38]
  wire  _new_s_T = ~adder_io_out_c_reg_0; // @[FloatingPointDesigns.scala 1501:15]
  wire  new_s = ~adder_io_out_c_reg_0 & (sign_reg_5_0 | sign_reg_5_1) | sign_reg_5_0 & sign_reg_5_1; // @[FloatingPointDesigns.scala 1501:75]
  wire  _D_T_1 = sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1508:53]
  wire  D = _new_s_T | sign_reg_5_0 ^ sign_reg_5_1; // @[FloatingPointDesigns.scala 1508:35]
  wire  E = _new_s_T & ~adder_io_out_s_reg_0[23] | _new_s_T & ~_D_T_1 | adder_io_out_c_reg_0 & adder_io_out_s_reg_0[23]
     & _D_T_1; // @[FloatingPointDesigns.scala 1510:134]
  reg [23:0] cmpl_adder_io_out_s_reg_0; // @[FloatingPointDesigns.scala 1512:42]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T = ~adder_io_out_s_reg_1; // @[FloatingPointDesigns.scala 1515:43]
  wire [23:0] _cmpl_adder_io_out_s_reg_0_T_2 = 24'h1 + _cmpl_adder_io_out_s_reg_0_T; // @[FloatingPointDesigns.scala 1515:41]
  wire [1:0] _adder_result_T = {sign_reg_7_1,sign_reg_7_0}; // @[FloatingPointDesigns.scala 1519:53]
  wire [1:0] _leadingOne_T_25 = adder_result_reg_0[2] ? 2'h2 : {{1'd0}, adder_result_reg_0[1]}; // @[FloatingPointDesigns.scala 1522:70]
  wire [1:0] _leadingOne_T_26 = adder_result_reg_0[3] ? 2'h3 : _leadingOne_T_25; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_27 = adder_result_reg_0[4] ? 3'h4 : {{1'd0}, _leadingOne_T_26}; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_28 = adder_result_reg_0[5] ? 3'h5 : _leadingOne_T_27; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_29 = adder_result_reg_0[6] ? 3'h6 : _leadingOne_T_28; // @[FloatingPointDesigns.scala 1522:70]
  wire [2:0] _leadingOne_T_30 = adder_result_reg_0[7] ? 3'h7 : _leadingOne_T_29; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_31 = adder_result_reg_0[8] ? 4'h8 : {{1'd0}, _leadingOne_T_30}; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_32 = adder_result_reg_0[9] ? 4'h9 : _leadingOne_T_31; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_33 = adder_result_reg_0[10] ? 4'ha : _leadingOne_T_32; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_34 = adder_result_reg_0[11] ? 4'hb : _leadingOne_T_33; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_35 = adder_result_reg_0[12] ? 4'hc : _leadingOne_T_34; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_36 = adder_result_reg_0[13] ? 4'hd : _leadingOne_T_35; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_37 = adder_result_reg_0[14] ? 4'he : _leadingOne_T_36; // @[FloatingPointDesigns.scala 1522:70]
  wire [3:0] _leadingOne_T_38 = adder_result_reg_0[15] ? 4'hf : _leadingOne_T_37; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_39 = adder_result_reg_0[16] ? 5'h10 : {{1'd0}, _leadingOne_T_38}; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_40 = adder_result_reg_0[17] ? 5'h11 : _leadingOne_T_39; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_41 = adder_result_reg_0[18] ? 5'h12 : _leadingOne_T_40; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_42 = adder_result_reg_0[19] ? 5'h13 : _leadingOne_T_41; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_43 = adder_result_reg_0[20] ? 5'h14 : _leadingOne_T_42; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_44 = adder_result_reg_0[21] ? 5'h15 : _leadingOne_T_43; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_45 = adder_result_reg_0[22] ? 5'h16 : _leadingOne_T_44; // @[FloatingPointDesigns.scala 1522:70]
  wire [4:0] _leadingOne_T_46 = adder_result_reg_0[23] ? 5'h17 : _leadingOne_T_45; // @[FloatingPointDesigns.scala 1522:70]
  wire [5:0] leadingOne = _leadingOne_T_46 + 5'h1; // @[FloatingPointDesigns.scala 1522:77]
  wire [5:0] _subber2_io_in_b_T_1 = 6'h18 - leadingOne_reg_0; // @[FloatingPointDesigns.scala 1525:42]
  wire [7:0] exp_0 = _GEN_1[7:0]; // @[FloatingPointDesigns.scala 1387:19]
  wire [7:0] exp_1 = _GEN_3[7:0]; // @[FloatingPointDesigns.scala 1387:19]
  wire [7:0] _GEN_24 = subber_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1538:27 1419:35]
  wire  _GEN_25 = subber_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1539:27 1420:35]
  wire [23:0] _GEN_35 = adder_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1554:29 1429:37]
  wire  _GEN_36 = adder_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1555:29 1430:37]
  wire [7:0] _GEN_39 = subber2_io_out_s; // @[FloatingPointDesigns.scala 1529:19 1561:28 1445:36]
  wire  _GEN_40 = subber2_io_out_c; // @[FloatingPointDesigns.scala 1529:19 1562:28 1446:36]
  reg [31:0] reg_out_s; // @[FloatingPointDesigns.scala 1596:28]
  wire [8:0] _GEN_169 = {{1'd0}, ref_exp_reg_7}; // @[FloatingPointDesigns.scala 1613:29]
  wire [23:0] _new_out_frac_reg_0_T_2 = 24'h800000 - 24'h1; // @[FloatingPointDesigns.scala 1615:60]
  wire [7:0] _new_out_exp_reg_0_T_3 = ref_exp_reg_7 + 8'h1; // @[FloatingPointDesigns.scala 1617:48]
  wire [8:0] _GEN_142 = _GEN_169 == _T_2 ? _T_2 : {{1'd0}, _new_out_exp_reg_0_T_3}; // @[FloatingPointDesigns.scala 1613:66 1614:30 1617:30]
  wire [23:0] _GEN_143 = _GEN_169 == _T_2 ? _new_out_frac_reg_0_T_2 : {{1'd0}, adder_result_reg_2[23:1]}; // @[FloatingPointDesigns.scala 1613:66 1615:31 1618:31]
  wire [5:0] _new_out_frac_reg_0_T_6 = 6'h18 - leadingOne_reg_1; // @[FloatingPointDesigns.scala 1631:94]
  wire [85:0] _GEN_4 = {{63'd0}, adder_result_reg_2[22:0]}; // @[FloatingPointDesigns.scala 1631:73]
  wire [85:0] _new_out_frac_reg_0_T_7 = _GEN_4 << _new_out_frac_reg_0_T_6; // @[FloatingPointDesigns.scala 1631:73]
  wire [7:0] _GEN_144 = subber2_out_c_reg_0 ? 8'h1 : subber2_out_s_reg_0; // @[FloatingPointDesigns.scala 1626:46 1627:32 1630:32]
  wire [85:0] _GEN_145 = subber2_out_c_reg_0 ? 86'h0 : _new_out_frac_reg_0_T_7; // @[FloatingPointDesigns.scala 1626:46 1628:33 1631:33]
  wire [7:0] _GEN_146 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 8'h0 : _GEN_144; // @[FloatingPointDesigns.scala 1622:184 1623:30]
  wire [85:0] _GEN_147 = leadingOne_reg_1 == 6'h1 & adder_result_reg_2 == 24'h0 & ((sign_reg_10_0 ^ sign_reg_10_1) &
    io_in_a_reg_10[30:0] == io_in_b_reg_10[30:0]) ? 86'h0 : _GEN_145; // @[FloatingPointDesigns.scala 1622:184 1624:31]
  wire  _GEN_148 = D_reg_4 ? new_s_reg_4 : new_s_reg_5; // @[FloatingPointDesigns.scala 1620:36 1621:22 1432:35]
  wire [7:0] _GEN_149 = D_reg_4 ? _GEN_146 : new_out_exp_reg_0; // @[FloatingPointDesigns.scala 1434:35 1620:36]
  wire [85:0] _GEN_150 = D_reg_4 ? _GEN_147 : {{63'd0}, new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1433:35 1620:36]
  wire  _GEN_151 = ~D_reg_4 ? new_s_reg_4 : _GEN_148; // @[FloatingPointDesigns.scala 1611:36 1612:22]
  wire [8:0] _GEN_152 = ~D_reg_4 ? _GEN_142 : {{1'd0}, _GEN_149}; // @[FloatingPointDesigns.scala 1611:36]
  wire [85:0] _GEN_153 = ~D_reg_4 ? {{62'd0}, _GEN_143} : _GEN_150; // @[FloatingPointDesigns.scala 1611:36]
  wire [8:0] _GEN_155 = E_reg_4 ? {{1'd0}, ref_exp_reg_7} : _GEN_152; // @[FloatingPointDesigns.scala 1607:36 1609:28]
  wire [85:0] _GEN_156 = E_reg_4 ? {{63'd0}, adder_result_reg_2[22:0]} : _GEN_153; // @[FloatingPointDesigns.scala 1607:36 1610:29]
  wire [85:0] _GEN_158 = sub_exp_reg_7 >= 8'h17 ? {{63'd0}, ref_frac_reg_7} : _GEN_156; // @[FloatingPointDesigns.scala 1603:48 1605:29]
  wire [8:0] _GEN_159 = sub_exp_reg_7 >= 8'h17 ? {{1'd0}, ref_exp_reg_7} : _GEN_155; // @[FloatingPointDesigns.scala 1603:48 1606:28]
  wire [8:0] _GEN_161 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 9'h0 : _GEN_159; // @[FloatingPointDesigns.scala 1599:86 1601:28]
  wire [85:0] _GEN_162 = io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0 ? 86'h0 : _GEN_158; // @[FloatingPointDesigns.scala 1599:86 1602:29]
  wire [31:0] _reg_out_s_T_1 = {new_s_reg_5,new_out_exp_reg_0,new_out_frac_reg_0}; // @[FloatingPointDesigns.scala 1635:55]
  wire [85:0] _GEN_170 = reset ? 86'h0 : _GEN_162; // @[FloatingPointDesigns.scala 1433:{35,35}]
  wire [8:0] _GEN_171 = reset ? 9'h0 : _GEN_161; // @[FloatingPointDesigns.scala 1434:{35,35}]
  full_subber subber ( // @[FloatingPointDesigns.scala 1456:24]
    .io_in_a(subber_io_in_a),
    .io_in_b(subber_io_in_b),
    .io_out_s(subber_io_out_s),
    .io_out_c(subber_io_out_c)
  );
  full_adder_64 adder ( // @[FloatingPointDesigns.scala 1462:23]
    .io_in_a(adder_io_in_a),
    .io_in_b(adder_io_in_b),
    .io_out_s(adder_io_out_s),
    .io_out_c(adder_io_out_c)
  );
  full_subber subber2 ( // @[FloatingPointDesigns.scala 1523:25]
    .io_in_a(subber2_io_in_a),
    .io_in_b(subber2_io_in_b),
    .io_out_s(subber2_io_out_s),
    .io_out_c(subber2_io_out_c)
  );
  assign io_out_s = reg_out_s; // @[FloatingPointDesigns.scala 1597:14]
  assign subber_io_in_a = exp_reg_0_0; // @[FloatingPointDesigns.scala 1457:20]
  assign subber_io_in_b = exp_reg_0_1; // @[FloatingPointDesigns.scala 1458:20]
  assign adder_io_in_a = _adder_io_in_a_T == 2'h1 ? cmpl_wire_temp_add_in_reg_0_0 : wire_temp_add_in_reg_1_0; // @[FloatingPointDesigns.scala 1494:25]
  assign adder_io_in_b = _adder_io_in_a_T == 2'h2 ? cmpl_wire_temp_add_in_reg_0_1 : wire_temp_add_in_reg_1_1; // @[FloatingPointDesigns.scala 1495:25]
  assign subber2_io_in_a = ref_exp_reg_6; // @[FloatingPointDesigns.scala 1524:21]
  assign subber2_io_in_b = {{2'd0}, _subber2_io_in_b_T_1}; // @[FloatingPointDesigns.scala 1525:21]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_0_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_0_0 <= sign_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_0_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_0_1 <= sign_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_1_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_1_0 <= sign_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_1_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_1_1 <= sign_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_2_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_2_0 <= sign_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_2_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_2_1 <= sign_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_3_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_3_0 <= sign_reg_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_3_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_3_1 <= sign_reg_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_4_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_4_0 <= sign_reg_3_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_4_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_4_1 <= sign_reg_3_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_5_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_5_0 <= sign_reg_4_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_5_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_5_1 <= sign_reg_4_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_6_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_6_0 <= sign_reg_5_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_6_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_6_1 <= sign_reg_5_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_7_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_7_0 <= sign_reg_6_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_7_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_7_1 <= sign_reg_6_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_8_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_8_0 <= sign_reg_7_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_8_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_8_1 <= sign_reg_7_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_9_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_9_0 <= sign_reg_8_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_9_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_9_1 <= sign_reg_8_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_10_0 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_10_0 <= sign_reg_9_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1414:28]
      sign_reg_10_1 <= 1'h0; // @[FloatingPointDesigns.scala 1414:28]
    end else begin
      sign_reg_10_1 <= sign_reg_9_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_0_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_0_0 <= exp_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_0_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_0_1 <= exp_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_1_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_1_0 <= exp_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_1_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_1_1 <= exp_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_2_0 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_2_0 <= exp_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1415:28]
      exp_reg_2_1 <= 8'h0; // @[FloatingPointDesigns.scala 1415:28]
    end else begin
      exp_reg_2_1 <= exp_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_0_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_0_0 <= frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_0_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_0_1 <= frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_1_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_1_0 <= frac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_1_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_1_1 <= frac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_2_0 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_2_0 <= frac_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1416:28]
      frac_reg_2_1 <= 23'h0; // @[FloatingPointDesigns.scala 1416:28]
    end else begin
      frac_reg_2_1 <= frac_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_0_0 <= whole_frac_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_0_1 <= whole_frac_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_1_0 <= wfrac_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_1_1 <= wfrac_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_2_0 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_2_0 <= wfrac_reg_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1417:28]
      wfrac_reg_2_1 <= 24'h0; // @[FloatingPointDesigns.scala 1417:28]
    end else begin
      wfrac_reg_2_1 <= wfrac_reg_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1419:35]
      subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1419:35]
    end else begin
      subber_out_s_reg_0 <= _GEN_24;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1419:35]
      subber_out_s_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1419:35]
    end else begin
      subber_out_s_reg_1 <= subber_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1420:35]
      subber_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1420:35]
    end else begin
      subber_out_c_reg_0 <= _GEN_25;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1420:35]
      subber_out_c_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1420:35]
    end else begin
      subber_out_c_reg_1 <= subber_out_c_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      wire_temp_add_in_reg_0_0 <= _wire_temp_add_in_0_T; // @[FloatingPointDesigns.scala 1477:27]
    end else begin
      wire_temp_add_in_reg_0_0 <= wfrac_reg_2_0; // @[FloatingPointDesigns.scala 1484:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      wire_temp_add_in_reg_0_1 <= wfrac_reg_2_1; // @[FloatingPointDesigns.scala 1478:27]
    end else begin
      wire_temp_add_in_reg_0_1 <= _wire_temp_add_in_1_T; // @[FloatingPointDesigns.scala 1485:27]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_1_0 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else begin
      wire_temp_add_in_reg_1_0 <= wire_temp_add_in_reg_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1422:39]
      wire_temp_add_in_reg_1_1 <= 24'h0; // @[FloatingPointDesigns.scala 1422:39]
    end else begin
      wire_temp_add_in_reg_1_1 <= wire_temp_add_in_reg_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_s_reg_0 <= sign_reg_2_1; // @[FloatingPointDesigns.scala 1475:13]
    end else begin
      ref_s_reg_0 <= sign_reg_2_0; // @[FloatingPointDesigns.scala 1482:13]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_1 <= ref_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_2 <= ref_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_3 <= ref_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_4 <= ref_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_5 <= ref_s_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_6 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_6 <= ref_s_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1424:31]
      ref_s_reg_7 <= 1'h0; // @[FloatingPointDesigns.scala 1424:31]
    end else begin
      ref_s_reg_7 <= ref_s_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_0 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_frac_reg_0 <= frac_reg_2_1; // @[FloatingPointDesigns.scala 1476:16]
    end else begin
      ref_frac_reg_0 <= frac_reg_2_0; // @[FloatingPointDesigns.scala 1483:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_1 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_1 <= ref_frac_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_2 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_2 <= ref_frac_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_3 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_3 <= ref_frac_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_4 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_4 <= ref_frac_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_5 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_5 <= ref_frac_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_6 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_6 <= ref_frac_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1425:31]
      ref_frac_reg_7 <= 23'h0; // @[FloatingPointDesigns.scala 1425:31]
    end else begin
      ref_frac_reg_7 <= ref_frac_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      ref_exp_reg_0 <= exp_reg_2_1; // @[FloatingPointDesigns.scala 1473:15]
    end else begin
      ref_exp_reg_0 <= exp_reg_2_0; // @[FloatingPointDesigns.scala 1480:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_1 <= ref_exp_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_2 <= ref_exp_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_3 <= ref_exp_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_4 <= ref_exp_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_5 <= ref_exp_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_6 <= ref_exp_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1426:31]
      ref_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1426:31]
    end else begin
      ref_exp_reg_7 <= ref_exp_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else if (subber_out_c_reg_1) begin // @[FloatingPointDesigns.scala 1472:39]
      sub_exp_reg_0 <= cmpl_subber_out_s_reg_0; // @[FloatingPointDesigns.scala 1474:15]
    end else begin
      sub_exp_reg_0 <= subber_out_s_reg_1; // @[FloatingPointDesigns.scala 1481:15]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_1 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_1 <= sub_exp_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_2 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_2 <= sub_exp_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_3 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_3 <= sub_exp_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_4 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_4 <= sub_exp_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_5 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_5 <= sub_exp_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_6 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_6 <= sub_exp_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1427:31]
      sub_exp_reg_7 <= 8'h0; // @[FloatingPointDesigns.scala 1427:31]
    end else begin
      sub_exp_reg_7 <= sub_exp_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_0 <= _GEN_35;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_1 <= adder_io_out_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1429:37]
      adder_io_out_s_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1429:37]
    end else begin
      adder_io_out_s_reg_2 <= adder_io_out_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1430:37]
      adder_io_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1430:37]
    end else begin
      adder_io_out_c_reg_0 <= _GEN_36;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_0 <= new_s;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_1 <= new_s_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_2 <= new_s_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_3 <= new_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else begin
      new_s_reg_4 <= new_s_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1432:35]
      new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1432:35]
    end else if (io_in_a_reg_10[30:0] == 31'h0 & io_in_b_reg_10[30:0] == 31'h0) begin // @[FloatingPointDesigns.scala 1599:86]
      new_s_reg_5 <= 1'h0; // @[FloatingPointDesigns.scala 1600:22]
    end else if (sub_exp_reg_7 >= 8'h17) begin // @[FloatingPointDesigns.scala 1603:48]
      new_s_reg_5 <= ref_s_reg_7; // @[FloatingPointDesigns.scala 1604:22]
    end else if (E_reg_4) begin // @[FloatingPointDesigns.scala 1607:36]
      new_s_reg_5 <= new_s_reg_4; // @[FloatingPointDesigns.scala 1608:22]
    end else begin
      new_s_reg_5 <= _GEN_151;
    end
    new_out_frac_reg_0 <= _GEN_170[22:0]; // @[FloatingPointDesigns.scala 1433:{35,35}]
    new_out_exp_reg_0 <= _GEN_171[7:0]; // @[FloatingPointDesigns.scala 1434:{35,35}]
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_0 <= E;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_1 <= E_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_2 <= E_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_3 <= E_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1435:24]
      E_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1435:24]
    end else begin
      E_reg_4 <= E_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_0 <= D;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_1 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_1 <= D_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_2 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_2 <= D_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_3 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_3 <= D_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1436:24]
      D_reg_4 <= 1'h0; // @[FloatingPointDesigns.scala 1436:24]
    end else begin
      D_reg_4 <= D_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else if (new_s_reg_1 & ^_adder_result_T) begin // @[FloatingPointDesigns.scala 1519:24]
      adder_result_reg_0 <= cmpl_adder_io_out_s_reg_0;
    end else begin
      adder_result_reg_0 <= adder_io_out_s_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_1 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else begin
      adder_result_reg_1 <= adder_result_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1438:35]
      adder_result_reg_2 <= 24'h0; // @[FloatingPointDesigns.scala 1438:35]
    end else begin
      adder_result_reg_2 <= adder_result_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1440:33]
      leadingOne_reg_0 <= 6'h0; // @[FloatingPointDesigns.scala 1440:33]
    end else begin
      leadingOne_reg_0 <= leadingOne;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1440:33]
      leadingOne_reg_1 <= 6'h0; // @[FloatingPointDesigns.scala 1440:33]
    end else begin
      leadingOne_reg_1 <= leadingOne_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_0 <= io_in_a;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_1 <= io_in_a_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_2 <= io_in_a_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_3 <= io_in_a_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_4 <= io_in_a_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_5 <= io_in_a_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_6 <= io_in_a_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_7 <= io_in_a_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_8 <= io_in_a_reg_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_9 <= io_in_a_reg_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1442:30]
      io_in_a_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1442:30]
    end else begin
      io_in_a_reg_10 <= io_in_a_reg_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_0 <= io_in_b;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_1 <= io_in_b_reg_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_2 <= io_in_b_reg_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_3 <= io_in_b_reg_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_4 <= io_in_b_reg_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_5 <= io_in_b_reg_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_6 <= io_in_b_reg_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_7 <= io_in_b_reg_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_8 <= io_in_b_reg_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_9 <= io_in_b_reg_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1443:30]
      io_in_b_reg_10 <= 32'h0; // @[FloatingPointDesigns.scala 1443:30]
    end else begin
      io_in_b_reg_10 <= io_in_b_reg_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1445:36]
      subber2_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1445:36]
    end else begin
      subber2_out_s_reg_0 <= _GEN_39;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1446:36]
      subber2_out_c_reg_0 <= 1'h0; // @[FloatingPointDesigns.scala 1446:36]
    end else begin
      subber2_out_c_reg_0 <= _GEN_40;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1467:40]
      cmpl_subber_out_s_reg_0 <= 8'h0; // @[FloatingPointDesigns.scala 1467:40]
    end else begin
      cmpl_subber_out_s_reg_0 <= _cmpl_subber_out_s_reg_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1488:44]
      cmpl_wire_temp_add_in_reg_0_0 <= 24'h0; // @[FloatingPointDesigns.scala 1488:44]
    end else begin
      cmpl_wire_temp_add_in_reg_0_0 <= _cmpl_wire_temp_add_in_reg_0_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1488:44]
      cmpl_wire_temp_add_in_reg_0_1 <= 24'h0; // @[FloatingPointDesigns.scala 1488:44]
    end else begin
      cmpl_wire_temp_add_in_reg_0_1 <= _cmpl_wire_temp_add_in_reg_0_1_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1512:42]
      cmpl_adder_io_out_s_reg_0 <= 24'h0; // @[FloatingPointDesigns.scala 1512:42]
    end else begin
      cmpl_adder_io_out_s_reg_0 <= _cmpl_adder_io_out_s_reg_0_T_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1596:28]
      reg_out_s <= 32'h0; // @[FloatingPointDesigns.scala 1596:28]
    end else begin
      reg_out_s <= _reg_out_s_T_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  sign_reg_0_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  sign_reg_0_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  sign_reg_1_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  sign_reg_1_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  sign_reg_2_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  sign_reg_2_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  sign_reg_3_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  sign_reg_3_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  sign_reg_4_0 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  sign_reg_4_1 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  sign_reg_5_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  sign_reg_5_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  sign_reg_6_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  sign_reg_6_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  sign_reg_7_0 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  sign_reg_7_1 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  sign_reg_8_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  sign_reg_8_1 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sign_reg_9_0 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sign_reg_9_1 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  sign_reg_10_0 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  sign_reg_10_1 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  exp_reg_0_0 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  exp_reg_0_1 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  exp_reg_1_0 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  exp_reg_1_1 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  exp_reg_2_0 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  exp_reg_2_1 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  frac_reg_0_0 = _RAND_28[22:0];
  _RAND_29 = {1{`RANDOM}};
  frac_reg_0_1 = _RAND_29[22:0];
  _RAND_30 = {1{`RANDOM}};
  frac_reg_1_0 = _RAND_30[22:0];
  _RAND_31 = {1{`RANDOM}};
  frac_reg_1_1 = _RAND_31[22:0];
  _RAND_32 = {1{`RANDOM}};
  frac_reg_2_0 = _RAND_32[22:0];
  _RAND_33 = {1{`RANDOM}};
  frac_reg_2_1 = _RAND_33[22:0];
  _RAND_34 = {1{`RANDOM}};
  wfrac_reg_0_0 = _RAND_34[23:0];
  _RAND_35 = {1{`RANDOM}};
  wfrac_reg_0_1 = _RAND_35[23:0];
  _RAND_36 = {1{`RANDOM}};
  wfrac_reg_1_0 = _RAND_36[23:0];
  _RAND_37 = {1{`RANDOM}};
  wfrac_reg_1_1 = _RAND_37[23:0];
  _RAND_38 = {1{`RANDOM}};
  wfrac_reg_2_0 = _RAND_38[23:0];
  _RAND_39 = {1{`RANDOM}};
  wfrac_reg_2_1 = _RAND_39[23:0];
  _RAND_40 = {1{`RANDOM}};
  subber_out_s_reg_0 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  subber_out_s_reg_1 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  subber_out_c_reg_0 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  subber_out_c_reg_1 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_0 = _RAND_44[23:0];
  _RAND_45 = {1{`RANDOM}};
  wire_temp_add_in_reg_0_1 = _RAND_45[23:0];
  _RAND_46 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_0 = _RAND_46[23:0];
  _RAND_47 = {1{`RANDOM}};
  wire_temp_add_in_reg_1_1 = _RAND_47[23:0];
  _RAND_48 = {1{`RANDOM}};
  ref_s_reg_0 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  ref_s_reg_1 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  ref_s_reg_2 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  ref_s_reg_3 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  ref_s_reg_4 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  ref_s_reg_5 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  ref_s_reg_6 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  ref_s_reg_7 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  ref_frac_reg_0 = _RAND_56[22:0];
  _RAND_57 = {1{`RANDOM}};
  ref_frac_reg_1 = _RAND_57[22:0];
  _RAND_58 = {1{`RANDOM}};
  ref_frac_reg_2 = _RAND_58[22:0];
  _RAND_59 = {1{`RANDOM}};
  ref_frac_reg_3 = _RAND_59[22:0];
  _RAND_60 = {1{`RANDOM}};
  ref_frac_reg_4 = _RAND_60[22:0];
  _RAND_61 = {1{`RANDOM}};
  ref_frac_reg_5 = _RAND_61[22:0];
  _RAND_62 = {1{`RANDOM}};
  ref_frac_reg_6 = _RAND_62[22:0];
  _RAND_63 = {1{`RANDOM}};
  ref_frac_reg_7 = _RAND_63[22:0];
  _RAND_64 = {1{`RANDOM}};
  ref_exp_reg_0 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  ref_exp_reg_1 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  ref_exp_reg_2 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  ref_exp_reg_3 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  ref_exp_reg_4 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  ref_exp_reg_5 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  ref_exp_reg_6 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  ref_exp_reg_7 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  sub_exp_reg_0 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  sub_exp_reg_1 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  sub_exp_reg_2 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  sub_exp_reg_3 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  sub_exp_reg_4 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  sub_exp_reg_5 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  sub_exp_reg_6 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  sub_exp_reg_7 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  adder_io_out_s_reg_0 = _RAND_80[23:0];
  _RAND_81 = {1{`RANDOM}};
  adder_io_out_s_reg_1 = _RAND_81[23:0];
  _RAND_82 = {1{`RANDOM}};
  adder_io_out_s_reg_2 = _RAND_82[23:0];
  _RAND_83 = {1{`RANDOM}};
  adder_io_out_c_reg_0 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  new_s_reg_0 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  new_s_reg_1 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  new_s_reg_2 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  new_s_reg_3 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  new_s_reg_4 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  new_s_reg_5 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  new_out_frac_reg_0 = _RAND_90[22:0];
  _RAND_91 = {1{`RANDOM}};
  new_out_exp_reg_0 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  E_reg_0 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  E_reg_1 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  E_reg_2 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  E_reg_3 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  E_reg_4 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  D_reg_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  D_reg_1 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  D_reg_2 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  D_reg_3 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  D_reg_4 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  adder_result_reg_0 = _RAND_102[23:0];
  _RAND_103 = {1{`RANDOM}};
  adder_result_reg_1 = _RAND_103[23:0];
  _RAND_104 = {1{`RANDOM}};
  adder_result_reg_2 = _RAND_104[23:0];
  _RAND_105 = {1{`RANDOM}};
  leadingOne_reg_0 = _RAND_105[5:0];
  _RAND_106 = {1{`RANDOM}};
  leadingOne_reg_1 = _RAND_106[5:0];
  _RAND_107 = {1{`RANDOM}};
  io_in_a_reg_0 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  io_in_a_reg_1 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  io_in_a_reg_2 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  io_in_a_reg_3 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  io_in_a_reg_4 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  io_in_a_reg_5 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  io_in_a_reg_6 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  io_in_a_reg_7 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  io_in_a_reg_8 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  io_in_a_reg_9 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  io_in_a_reg_10 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  io_in_b_reg_0 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  io_in_b_reg_1 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  io_in_b_reg_2 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  io_in_b_reg_3 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  io_in_b_reg_4 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  io_in_b_reg_5 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  io_in_b_reg_6 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  io_in_b_reg_7 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  io_in_b_reg_8 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  io_in_b_reg_9 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  io_in_b_reg_10 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  subber2_out_s_reg_0 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  subber2_out_c_reg_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cmpl_subber_out_s_reg_0 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_0 = _RAND_132[23:0];
  _RAND_133 = {1{`RANDOM}};
  cmpl_wire_temp_add_in_reg_0_1 = _RAND_133[23:0];
  _RAND_134 = {1{`RANDOM}};
  cmpl_adder_io_out_s_reg_0 = _RAND_134[23:0];
  _RAND_135 = {1{`RANDOM}};
  reg_out_s = _RAND_135[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_DDOT_dp(
  input         clock,
  input         reset,
  input  [31:0] io_in_a_0,
  input  [31:0] io_in_a_1,
  input  [31:0] io_in_a_2,
  input  [31:0] io_in_a_3,
  input  [31:0] io_in_a_4,
  input  [31:0] io_in_a_5,
  input  [31:0] io_in_a_6,
  input  [31:0] io_in_a_7,
  input  [31:0] io_in_a_8,
  input  [31:0] io_in_a_9,
  input  [31:0] io_in_a_10,
  input  [31:0] io_in_a_11,
  input  [31:0] io_in_a_12,
  input  [31:0] io_in_a_13,
  input  [31:0] io_in_a_14,
  input  [31:0] io_in_a_15,
  input  [31:0] io_in_a_16,
  input  [31:0] io_in_a_17,
  input  [31:0] io_in_a_18,
  input  [31:0] io_in_a_19,
  input  [31:0] io_in_a_20,
  input  [31:0] io_in_a_21,
  input  [31:0] io_in_a_22,
  input  [31:0] io_in_a_23,
  input  [31:0] io_in_a_24,
  input  [31:0] io_in_a_25,
  input  [31:0] io_in_a_26,
  input  [31:0] io_in_a_27,
  input  [31:0] io_in_a_28,
  input  [31:0] io_in_a_29,
  input  [31:0] io_in_a_30,
  input  [31:0] io_in_a_31,
  input  [31:0] io_in_a_32,
  input  [31:0] io_in_a_33,
  input  [31:0] io_in_a_34,
  input  [31:0] io_in_a_35,
  input  [31:0] io_in_a_36,
  input  [31:0] io_in_a_37,
  input  [31:0] io_in_a_38,
  input  [31:0] io_in_a_39,
  input  [31:0] io_in_a_40,
  input  [31:0] io_in_a_41,
  input  [31:0] io_in_a_42,
  input  [31:0] io_in_a_43,
  input  [31:0] io_in_a_44,
  input  [31:0] io_in_a_45,
  input  [31:0] io_in_a_46,
  input  [31:0] io_in_a_47,
  input  [31:0] io_in_a_48,
  input  [31:0] io_in_a_49,
  input  [31:0] io_in_a_50,
  input  [31:0] io_in_a_51,
  input  [31:0] io_in_a_52,
  input  [31:0] io_in_a_53,
  input  [31:0] io_in_a_54,
  input  [31:0] io_in_a_55,
  input  [31:0] io_in_a_56,
  input  [31:0] io_in_a_57,
  input  [31:0] io_in_a_58,
  input  [31:0] io_in_a_59,
  input  [31:0] io_in_a_60,
  input  [31:0] io_in_a_61,
  input  [31:0] io_in_a_62,
  input  [31:0] io_in_a_63,
  input  [31:0] io_in_b_0,
  input  [31:0] io_in_b_1,
  input  [31:0] io_in_b_2,
  input  [31:0] io_in_b_3,
  input  [31:0] io_in_b_4,
  input  [31:0] io_in_b_5,
  input  [31:0] io_in_b_6,
  input  [31:0] io_in_b_7,
  input  [31:0] io_in_b_8,
  input  [31:0] io_in_b_9,
  input  [31:0] io_in_b_10,
  input  [31:0] io_in_b_11,
  input  [31:0] io_in_b_12,
  input  [31:0] io_in_b_13,
  input  [31:0] io_in_b_14,
  input  [31:0] io_in_b_15,
  input  [31:0] io_in_b_16,
  input  [31:0] io_in_b_17,
  input  [31:0] io_in_b_18,
  input  [31:0] io_in_b_19,
  input  [31:0] io_in_b_20,
  input  [31:0] io_in_b_21,
  input  [31:0] io_in_b_22,
  input  [31:0] io_in_b_23,
  input  [31:0] io_in_b_24,
  input  [31:0] io_in_b_25,
  input  [31:0] io_in_b_26,
  input  [31:0] io_in_b_27,
  input  [31:0] io_in_b_28,
  input  [31:0] io_in_b_29,
  input  [31:0] io_in_b_30,
  input  [31:0] io_in_b_31,
  input  [31:0] io_in_b_32,
  input  [31:0] io_in_b_33,
  input  [31:0] io_in_b_34,
  input  [31:0] io_in_b_35,
  input  [31:0] io_in_b_36,
  input  [31:0] io_in_b_37,
  input  [31:0] io_in_b_38,
  input  [31:0] io_in_b_39,
  input  [31:0] io_in_b_40,
  input  [31:0] io_in_b_41,
  input  [31:0] io_in_b_42,
  input  [31:0] io_in_b_43,
  input  [31:0] io_in_b_44,
  input  [31:0] io_in_b_45,
  input  [31:0] io_in_b_46,
  input  [31:0] io_in_b_47,
  input  [31:0] io_in_b_48,
  input  [31:0] io_in_b_49,
  input  [31:0] io_in_b_50,
  input  [31:0] io_in_b_51,
  input  [31:0] io_in_b_52,
  input  [31:0] io_in_b_53,
  input  [31:0] io_in_b_54,
  input  [31:0] io_in_b_55,
  input  [31:0] io_in_b_56,
  input  [31:0] io_in_b_57,
  input  [31:0] io_in_b_58,
  input  [31:0] io_in_b_59,
  input  [31:0] io_in_b_60,
  input  [31:0] io_in_b_61,
  input  [31:0] io_in_b_62,
  input  [31:0] io_in_b_63,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_48_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_48_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_49_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_49_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_50_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_50_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_51_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_51_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_52_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_52_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_53_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_53_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_54_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_54_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_55_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_55_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_56_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_56_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_57_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_57_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_58_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_58_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_59_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_59_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_60_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_60_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_61_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_61_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_62_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_62_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_63_clock; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_multiplier_10ccs_63_reset; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2411:44]
  wire [31:0] FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2411:44]
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_1_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_1_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_2_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_2_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_3_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_3_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_4_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_4_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_5_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_5_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_6_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_6_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_7_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_7_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_8_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_8_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_9_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_9_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_10_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_10_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_11_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_11_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_12_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_12_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_13_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_13_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_14_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_14_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_15_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_15_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_16_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_16_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_17_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_17_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_18_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_18_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_19_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_19_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_20_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_20_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_21_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_21_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_22_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_22_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_23_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_23_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_24_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_24_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_25_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_25_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_26_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_26_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_27_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_27_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_28_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_28_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_29_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_29_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_30_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_30_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_31_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_31_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_32_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_32_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_33_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_33_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_34_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_34_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_35_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_35_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_36_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_36_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_37_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_37_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_38_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_38_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_39_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_39_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_40_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_40_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_41_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_41_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_42_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_42_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_43_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_43_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_44_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_44_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_45_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_45_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_46_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_46_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_47_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_47_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_48_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_48_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_49_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_49_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_50_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_50_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_51_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_51_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_52_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_52_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_53_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_53_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_54_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_54_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_55_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_55_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_56_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_56_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_57_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_57_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_58_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_58_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_59_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_59_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_60_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_60_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_61_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_61_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_62_clock; // @[FloatingPointDesigns.scala 2419:17]
  wire  FP_adder_13ccs_62_reset; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2419:17]
  wire [31:0] FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2419:17]
  reg [31:0] io_out_s_REG; // @[FloatingPointDesigns.scala 2468:26]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_48 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_48_clock),
    .reset(FP_multiplier_10ccs_48_reset),
    .io_in_a(FP_multiplier_10ccs_48_io_in_a),
    .io_in_b(FP_multiplier_10ccs_48_io_in_b),
    .io_out_s(FP_multiplier_10ccs_48_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_49 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_49_clock),
    .reset(FP_multiplier_10ccs_49_reset),
    .io_in_a(FP_multiplier_10ccs_49_io_in_a),
    .io_in_b(FP_multiplier_10ccs_49_io_in_b),
    .io_out_s(FP_multiplier_10ccs_49_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_50 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_50_clock),
    .reset(FP_multiplier_10ccs_50_reset),
    .io_in_a(FP_multiplier_10ccs_50_io_in_a),
    .io_in_b(FP_multiplier_10ccs_50_io_in_b),
    .io_out_s(FP_multiplier_10ccs_50_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_51 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_51_clock),
    .reset(FP_multiplier_10ccs_51_reset),
    .io_in_a(FP_multiplier_10ccs_51_io_in_a),
    .io_in_b(FP_multiplier_10ccs_51_io_in_b),
    .io_out_s(FP_multiplier_10ccs_51_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_52 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_52_clock),
    .reset(FP_multiplier_10ccs_52_reset),
    .io_in_a(FP_multiplier_10ccs_52_io_in_a),
    .io_in_b(FP_multiplier_10ccs_52_io_in_b),
    .io_out_s(FP_multiplier_10ccs_52_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_53 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_53_clock),
    .reset(FP_multiplier_10ccs_53_reset),
    .io_in_a(FP_multiplier_10ccs_53_io_in_a),
    .io_in_b(FP_multiplier_10ccs_53_io_in_b),
    .io_out_s(FP_multiplier_10ccs_53_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_54 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_54_clock),
    .reset(FP_multiplier_10ccs_54_reset),
    .io_in_a(FP_multiplier_10ccs_54_io_in_a),
    .io_in_b(FP_multiplier_10ccs_54_io_in_b),
    .io_out_s(FP_multiplier_10ccs_54_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_55 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_55_clock),
    .reset(FP_multiplier_10ccs_55_reset),
    .io_in_a(FP_multiplier_10ccs_55_io_in_a),
    .io_in_b(FP_multiplier_10ccs_55_io_in_b),
    .io_out_s(FP_multiplier_10ccs_55_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_56 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_56_clock),
    .reset(FP_multiplier_10ccs_56_reset),
    .io_in_a(FP_multiplier_10ccs_56_io_in_a),
    .io_in_b(FP_multiplier_10ccs_56_io_in_b),
    .io_out_s(FP_multiplier_10ccs_56_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_57 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_57_clock),
    .reset(FP_multiplier_10ccs_57_reset),
    .io_in_a(FP_multiplier_10ccs_57_io_in_a),
    .io_in_b(FP_multiplier_10ccs_57_io_in_b),
    .io_out_s(FP_multiplier_10ccs_57_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_58 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_58_clock),
    .reset(FP_multiplier_10ccs_58_reset),
    .io_in_a(FP_multiplier_10ccs_58_io_in_a),
    .io_in_b(FP_multiplier_10ccs_58_io_in_b),
    .io_out_s(FP_multiplier_10ccs_58_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_59 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_59_clock),
    .reset(FP_multiplier_10ccs_59_reset),
    .io_in_a(FP_multiplier_10ccs_59_io_in_a),
    .io_in_b(FP_multiplier_10ccs_59_io_in_b),
    .io_out_s(FP_multiplier_10ccs_59_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_60 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_60_clock),
    .reset(FP_multiplier_10ccs_60_reset),
    .io_in_a(FP_multiplier_10ccs_60_io_in_a),
    .io_in_b(FP_multiplier_10ccs_60_io_in_b),
    .io_out_s(FP_multiplier_10ccs_60_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_61 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_61_clock),
    .reset(FP_multiplier_10ccs_61_reset),
    .io_in_a(FP_multiplier_10ccs_61_io_in_a),
    .io_in_b(FP_multiplier_10ccs_61_io_in_b),
    .io_out_s(FP_multiplier_10ccs_61_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_62 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_62_clock),
    .reset(FP_multiplier_10ccs_62_reset),
    .io_in_a(FP_multiplier_10ccs_62_io_in_a),
    .io_in_b(FP_multiplier_10ccs_62_io_in_b),
    .io_out_s(FP_multiplier_10ccs_62_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_63 ( // @[FloatingPointDesigns.scala 2411:44]
    .clock(FP_multiplier_10ccs_63_clock),
    .reset(FP_multiplier_10ccs_63_reset),
    .io_in_a(FP_multiplier_10ccs_63_io_in_a),
    .io_in_b(FP_multiplier_10ccs_63_io_in_b),
    .io_out_s(FP_multiplier_10ccs_63_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_1 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_1_clock),
    .reset(FP_adder_13ccs_1_reset),
    .io_in_a(FP_adder_13ccs_1_io_in_a),
    .io_in_b(FP_adder_13ccs_1_io_in_b),
    .io_out_s(FP_adder_13ccs_1_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_2 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_2_clock),
    .reset(FP_adder_13ccs_2_reset),
    .io_in_a(FP_adder_13ccs_2_io_in_a),
    .io_in_b(FP_adder_13ccs_2_io_in_b),
    .io_out_s(FP_adder_13ccs_2_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_3 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_3_clock),
    .reset(FP_adder_13ccs_3_reset),
    .io_in_a(FP_adder_13ccs_3_io_in_a),
    .io_in_b(FP_adder_13ccs_3_io_in_b),
    .io_out_s(FP_adder_13ccs_3_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_4 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_4_clock),
    .reset(FP_adder_13ccs_4_reset),
    .io_in_a(FP_adder_13ccs_4_io_in_a),
    .io_in_b(FP_adder_13ccs_4_io_in_b),
    .io_out_s(FP_adder_13ccs_4_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_5 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_5_clock),
    .reset(FP_adder_13ccs_5_reset),
    .io_in_a(FP_adder_13ccs_5_io_in_a),
    .io_in_b(FP_adder_13ccs_5_io_in_b),
    .io_out_s(FP_adder_13ccs_5_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_6 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_6_clock),
    .reset(FP_adder_13ccs_6_reset),
    .io_in_a(FP_adder_13ccs_6_io_in_a),
    .io_in_b(FP_adder_13ccs_6_io_in_b),
    .io_out_s(FP_adder_13ccs_6_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_7 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_7_clock),
    .reset(FP_adder_13ccs_7_reset),
    .io_in_a(FP_adder_13ccs_7_io_in_a),
    .io_in_b(FP_adder_13ccs_7_io_in_b),
    .io_out_s(FP_adder_13ccs_7_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_8 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_8_clock),
    .reset(FP_adder_13ccs_8_reset),
    .io_in_a(FP_adder_13ccs_8_io_in_a),
    .io_in_b(FP_adder_13ccs_8_io_in_b),
    .io_out_s(FP_adder_13ccs_8_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_9 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_9_clock),
    .reset(FP_adder_13ccs_9_reset),
    .io_in_a(FP_adder_13ccs_9_io_in_a),
    .io_in_b(FP_adder_13ccs_9_io_in_b),
    .io_out_s(FP_adder_13ccs_9_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_10 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_10_clock),
    .reset(FP_adder_13ccs_10_reset),
    .io_in_a(FP_adder_13ccs_10_io_in_a),
    .io_in_b(FP_adder_13ccs_10_io_in_b),
    .io_out_s(FP_adder_13ccs_10_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_11 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_11_clock),
    .reset(FP_adder_13ccs_11_reset),
    .io_in_a(FP_adder_13ccs_11_io_in_a),
    .io_in_b(FP_adder_13ccs_11_io_in_b),
    .io_out_s(FP_adder_13ccs_11_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_12 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_12_clock),
    .reset(FP_adder_13ccs_12_reset),
    .io_in_a(FP_adder_13ccs_12_io_in_a),
    .io_in_b(FP_adder_13ccs_12_io_in_b),
    .io_out_s(FP_adder_13ccs_12_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_13 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_13_clock),
    .reset(FP_adder_13ccs_13_reset),
    .io_in_a(FP_adder_13ccs_13_io_in_a),
    .io_in_b(FP_adder_13ccs_13_io_in_b),
    .io_out_s(FP_adder_13ccs_13_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_14 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_14_clock),
    .reset(FP_adder_13ccs_14_reset),
    .io_in_a(FP_adder_13ccs_14_io_in_a),
    .io_in_b(FP_adder_13ccs_14_io_in_b),
    .io_out_s(FP_adder_13ccs_14_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_15 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_15_clock),
    .reset(FP_adder_13ccs_15_reset),
    .io_in_a(FP_adder_13ccs_15_io_in_a),
    .io_in_b(FP_adder_13ccs_15_io_in_b),
    .io_out_s(FP_adder_13ccs_15_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_16 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_16_clock),
    .reset(FP_adder_13ccs_16_reset),
    .io_in_a(FP_adder_13ccs_16_io_in_a),
    .io_in_b(FP_adder_13ccs_16_io_in_b),
    .io_out_s(FP_adder_13ccs_16_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_17 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_17_clock),
    .reset(FP_adder_13ccs_17_reset),
    .io_in_a(FP_adder_13ccs_17_io_in_a),
    .io_in_b(FP_adder_13ccs_17_io_in_b),
    .io_out_s(FP_adder_13ccs_17_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_18 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_18_clock),
    .reset(FP_adder_13ccs_18_reset),
    .io_in_a(FP_adder_13ccs_18_io_in_a),
    .io_in_b(FP_adder_13ccs_18_io_in_b),
    .io_out_s(FP_adder_13ccs_18_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_19 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_19_clock),
    .reset(FP_adder_13ccs_19_reset),
    .io_in_a(FP_adder_13ccs_19_io_in_a),
    .io_in_b(FP_adder_13ccs_19_io_in_b),
    .io_out_s(FP_adder_13ccs_19_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_20 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_20_clock),
    .reset(FP_adder_13ccs_20_reset),
    .io_in_a(FP_adder_13ccs_20_io_in_a),
    .io_in_b(FP_adder_13ccs_20_io_in_b),
    .io_out_s(FP_adder_13ccs_20_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_21 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_21_clock),
    .reset(FP_adder_13ccs_21_reset),
    .io_in_a(FP_adder_13ccs_21_io_in_a),
    .io_in_b(FP_adder_13ccs_21_io_in_b),
    .io_out_s(FP_adder_13ccs_21_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_22 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_22_clock),
    .reset(FP_adder_13ccs_22_reset),
    .io_in_a(FP_adder_13ccs_22_io_in_a),
    .io_in_b(FP_adder_13ccs_22_io_in_b),
    .io_out_s(FP_adder_13ccs_22_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_23 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_23_clock),
    .reset(FP_adder_13ccs_23_reset),
    .io_in_a(FP_adder_13ccs_23_io_in_a),
    .io_in_b(FP_adder_13ccs_23_io_in_b),
    .io_out_s(FP_adder_13ccs_23_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_24 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_24_clock),
    .reset(FP_adder_13ccs_24_reset),
    .io_in_a(FP_adder_13ccs_24_io_in_a),
    .io_in_b(FP_adder_13ccs_24_io_in_b),
    .io_out_s(FP_adder_13ccs_24_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_25 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_25_clock),
    .reset(FP_adder_13ccs_25_reset),
    .io_in_a(FP_adder_13ccs_25_io_in_a),
    .io_in_b(FP_adder_13ccs_25_io_in_b),
    .io_out_s(FP_adder_13ccs_25_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_26 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_26_clock),
    .reset(FP_adder_13ccs_26_reset),
    .io_in_a(FP_adder_13ccs_26_io_in_a),
    .io_in_b(FP_adder_13ccs_26_io_in_b),
    .io_out_s(FP_adder_13ccs_26_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_27 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_27_clock),
    .reset(FP_adder_13ccs_27_reset),
    .io_in_a(FP_adder_13ccs_27_io_in_a),
    .io_in_b(FP_adder_13ccs_27_io_in_b),
    .io_out_s(FP_adder_13ccs_27_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_28 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_28_clock),
    .reset(FP_adder_13ccs_28_reset),
    .io_in_a(FP_adder_13ccs_28_io_in_a),
    .io_in_b(FP_adder_13ccs_28_io_in_b),
    .io_out_s(FP_adder_13ccs_28_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_29 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_29_clock),
    .reset(FP_adder_13ccs_29_reset),
    .io_in_a(FP_adder_13ccs_29_io_in_a),
    .io_in_b(FP_adder_13ccs_29_io_in_b),
    .io_out_s(FP_adder_13ccs_29_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_30 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_30_clock),
    .reset(FP_adder_13ccs_30_reset),
    .io_in_a(FP_adder_13ccs_30_io_in_a),
    .io_in_b(FP_adder_13ccs_30_io_in_b),
    .io_out_s(FP_adder_13ccs_30_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_31 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_31_clock),
    .reset(FP_adder_13ccs_31_reset),
    .io_in_a(FP_adder_13ccs_31_io_in_a),
    .io_in_b(FP_adder_13ccs_31_io_in_b),
    .io_out_s(FP_adder_13ccs_31_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_32 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_32_clock),
    .reset(FP_adder_13ccs_32_reset),
    .io_in_a(FP_adder_13ccs_32_io_in_a),
    .io_in_b(FP_adder_13ccs_32_io_in_b),
    .io_out_s(FP_adder_13ccs_32_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_33 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_33_clock),
    .reset(FP_adder_13ccs_33_reset),
    .io_in_a(FP_adder_13ccs_33_io_in_a),
    .io_in_b(FP_adder_13ccs_33_io_in_b),
    .io_out_s(FP_adder_13ccs_33_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_34 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_34_clock),
    .reset(FP_adder_13ccs_34_reset),
    .io_in_a(FP_adder_13ccs_34_io_in_a),
    .io_in_b(FP_adder_13ccs_34_io_in_b),
    .io_out_s(FP_adder_13ccs_34_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_35 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_35_clock),
    .reset(FP_adder_13ccs_35_reset),
    .io_in_a(FP_adder_13ccs_35_io_in_a),
    .io_in_b(FP_adder_13ccs_35_io_in_b),
    .io_out_s(FP_adder_13ccs_35_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_36 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_36_clock),
    .reset(FP_adder_13ccs_36_reset),
    .io_in_a(FP_adder_13ccs_36_io_in_a),
    .io_in_b(FP_adder_13ccs_36_io_in_b),
    .io_out_s(FP_adder_13ccs_36_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_37 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_37_clock),
    .reset(FP_adder_13ccs_37_reset),
    .io_in_a(FP_adder_13ccs_37_io_in_a),
    .io_in_b(FP_adder_13ccs_37_io_in_b),
    .io_out_s(FP_adder_13ccs_37_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_38 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_38_clock),
    .reset(FP_adder_13ccs_38_reset),
    .io_in_a(FP_adder_13ccs_38_io_in_a),
    .io_in_b(FP_adder_13ccs_38_io_in_b),
    .io_out_s(FP_adder_13ccs_38_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_39 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_39_clock),
    .reset(FP_adder_13ccs_39_reset),
    .io_in_a(FP_adder_13ccs_39_io_in_a),
    .io_in_b(FP_adder_13ccs_39_io_in_b),
    .io_out_s(FP_adder_13ccs_39_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_40 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_40_clock),
    .reset(FP_adder_13ccs_40_reset),
    .io_in_a(FP_adder_13ccs_40_io_in_a),
    .io_in_b(FP_adder_13ccs_40_io_in_b),
    .io_out_s(FP_adder_13ccs_40_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_41 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_41_clock),
    .reset(FP_adder_13ccs_41_reset),
    .io_in_a(FP_adder_13ccs_41_io_in_a),
    .io_in_b(FP_adder_13ccs_41_io_in_b),
    .io_out_s(FP_adder_13ccs_41_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_42 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_42_clock),
    .reset(FP_adder_13ccs_42_reset),
    .io_in_a(FP_adder_13ccs_42_io_in_a),
    .io_in_b(FP_adder_13ccs_42_io_in_b),
    .io_out_s(FP_adder_13ccs_42_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_43 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_43_clock),
    .reset(FP_adder_13ccs_43_reset),
    .io_in_a(FP_adder_13ccs_43_io_in_a),
    .io_in_b(FP_adder_13ccs_43_io_in_b),
    .io_out_s(FP_adder_13ccs_43_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_44 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_44_clock),
    .reset(FP_adder_13ccs_44_reset),
    .io_in_a(FP_adder_13ccs_44_io_in_a),
    .io_in_b(FP_adder_13ccs_44_io_in_b),
    .io_out_s(FP_adder_13ccs_44_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_45 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_45_clock),
    .reset(FP_adder_13ccs_45_reset),
    .io_in_a(FP_adder_13ccs_45_io_in_a),
    .io_in_b(FP_adder_13ccs_45_io_in_b),
    .io_out_s(FP_adder_13ccs_45_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_46 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_46_clock),
    .reset(FP_adder_13ccs_46_reset),
    .io_in_a(FP_adder_13ccs_46_io_in_a),
    .io_in_b(FP_adder_13ccs_46_io_in_b),
    .io_out_s(FP_adder_13ccs_46_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_47 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_47_clock),
    .reset(FP_adder_13ccs_47_reset),
    .io_in_a(FP_adder_13ccs_47_io_in_a),
    .io_in_b(FP_adder_13ccs_47_io_in_b),
    .io_out_s(FP_adder_13ccs_47_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_48 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_48_clock),
    .reset(FP_adder_13ccs_48_reset),
    .io_in_a(FP_adder_13ccs_48_io_in_a),
    .io_in_b(FP_adder_13ccs_48_io_in_b),
    .io_out_s(FP_adder_13ccs_48_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_49 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_49_clock),
    .reset(FP_adder_13ccs_49_reset),
    .io_in_a(FP_adder_13ccs_49_io_in_a),
    .io_in_b(FP_adder_13ccs_49_io_in_b),
    .io_out_s(FP_adder_13ccs_49_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_50 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_50_clock),
    .reset(FP_adder_13ccs_50_reset),
    .io_in_a(FP_adder_13ccs_50_io_in_a),
    .io_in_b(FP_adder_13ccs_50_io_in_b),
    .io_out_s(FP_adder_13ccs_50_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_51 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_51_clock),
    .reset(FP_adder_13ccs_51_reset),
    .io_in_a(FP_adder_13ccs_51_io_in_a),
    .io_in_b(FP_adder_13ccs_51_io_in_b),
    .io_out_s(FP_adder_13ccs_51_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_52 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_52_clock),
    .reset(FP_adder_13ccs_52_reset),
    .io_in_a(FP_adder_13ccs_52_io_in_a),
    .io_in_b(FP_adder_13ccs_52_io_in_b),
    .io_out_s(FP_adder_13ccs_52_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_53 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_53_clock),
    .reset(FP_adder_13ccs_53_reset),
    .io_in_a(FP_adder_13ccs_53_io_in_a),
    .io_in_b(FP_adder_13ccs_53_io_in_b),
    .io_out_s(FP_adder_13ccs_53_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_54 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_54_clock),
    .reset(FP_adder_13ccs_54_reset),
    .io_in_a(FP_adder_13ccs_54_io_in_a),
    .io_in_b(FP_adder_13ccs_54_io_in_b),
    .io_out_s(FP_adder_13ccs_54_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_55 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_55_clock),
    .reset(FP_adder_13ccs_55_reset),
    .io_in_a(FP_adder_13ccs_55_io_in_a),
    .io_in_b(FP_adder_13ccs_55_io_in_b),
    .io_out_s(FP_adder_13ccs_55_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_56 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_56_clock),
    .reset(FP_adder_13ccs_56_reset),
    .io_in_a(FP_adder_13ccs_56_io_in_a),
    .io_in_b(FP_adder_13ccs_56_io_in_b),
    .io_out_s(FP_adder_13ccs_56_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_57 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_57_clock),
    .reset(FP_adder_13ccs_57_reset),
    .io_in_a(FP_adder_13ccs_57_io_in_a),
    .io_in_b(FP_adder_13ccs_57_io_in_b),
    .io_out_s(FP_adder_13ccs_57_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_58 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_58_clock),
    .reset(FP_adder_13ccs_58_reset),
    .io_in_a(FP_adder_13ccs_58_io_in_a),
    .io_in_b(FP_adder_13ccs_58_io_in_b),
    .io_out_s(FP_adder_13ccs_58_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_59 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_59_clock),
    .reset(FP_adder_13ccs_59_reset),
    .io_in_a(FP_adder_13ccs_59_io_in_a),
    .io_in_b(FP_adder_13ccs_59_io_in_b),
    .io_out_s(FP_adder_13ccs_59_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_60 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_60_clock),
    .reset(FP_adder_13ccs_60_reset),
    .io_in_a(FP_adder_13ccs_60_io_in_a),
    .io_in_b(FP_adder_13ccs_60_io_in_b),
    .io_out_s(FP_adder_13ccs_60_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_61 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_61_clock),
    .reset(FP_adder_13ccs_61_reset),
    .io_in_a(FP_adder_13ccs_61_io_in_a),
    .io_in_b(FP_adder_13ccs_61_io_in_b),
    .io_out_s(FP_adder_13ccs_61_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_62 ( // @[FloatingPointDesigns.scala 2419:17]
    .clock(FP_adder_13ccs_62_clock),
    .reset(FP_adder_13ccs_62_reset),
    .io_in_a(FP_adder_13ccs_62_io_in_a),
    .io_in_b(FP_adder_13ccs_62_io_in_b),
    .io_out_s(FP_adder_13ccs_62_io_out_s)
  );
  assign io_out_s = io_out_s_REG; // @[FloatingPointDesigns.scala 2468:16]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = io_in_a_0; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_io_in_b = io_in_b_0; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = io_in_a_1; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_1_io_in_b = io_in_b_1; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = io_in_a_2; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_2_io_in_b = io_in_b_2; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = io_in_a_3; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_3_io_in_b = io_in_b_3; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = io_in_a_4; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_4_io_in_b = io_in_b_4; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = io_in_a_5; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_5_io_in_b = io_in_b_5; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = io_in_a_6; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_6_io_in_b = io_in_b_6; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = io_in_a_7; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_7_io_in_b = io_in_b_7; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = io_in_a_8; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_8_io_in_b = io_in_b_8; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_a = io_in_a_9; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_9_io_in_b = io_in_b_9; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_a = io_in_a_10; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_10_io_in_b = io_in_b_10; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_a = io_in_a_11; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_11_io_in_b = io_in_b_11; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_a = io_in_a_12; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_12_io_in_b = io_in_b_12; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_a = io_in_a_13; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_13_io_in_b = io_in_b_13; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_a = io_in_a_14; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_14_io_in_b = io_in_b_14; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_a = io_in_a_15; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_15_io_in_b = io_in_b_15; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_a = io_in_a_16; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_16_io_in_b = io_in_b_16; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_a = io_in_a_17; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_17_io_in_b = io_in_b_17; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_a = io_in_a_18; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_18_io_in_b = io_in_b_18; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_a = io_in_a_19; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_19_io_in_b = io_in_b_19; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_a = io_in_a_20; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_20_io_in_b = io_in_b_20; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_a = io_in_a_21; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_21_io_in_b = io_in_b_21; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_a = io_in_a_22; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_22_io_in_b = io_in_b_22; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_a = io_in_a_23; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_23_io_in_b = io_in_b_23; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_a = io_in_a_24; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_24_io_in_b = io_in_b_24; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_a = io_in_a_25; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_25_io_in_b = io_in_b_25; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_a = io_in_a_26; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_26_io_in_b = io_in_b_26; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_a = io_in_a_27; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_27_io_in_b = io_in_b_27; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_a = io_in_a_28; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_28_io_in_b = io_in_b_28; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_a = io_in_a_29; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_29_io_in_b = io_in_b_29; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_a = io_in_a_30; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_30_io_in_b = io_in_b_30; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_a = io_in_a_31; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_31_io_in_b = io_in_b_31; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_a = io_in_a_32; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_32_io_in_b = io_in_b_32; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_a = io_in_a_33; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_33_io_in_b = io_in_b_33; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_a = io_in_a_34; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_34_io_in_b = io_in_b_34; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_a = io_in_a_35; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_35_io_in_b = io_in_b_35; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_a = io_in_a_36; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_36_io_in_b = io_in_b_36; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_a = io_in_a_37; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_37_io_in_b = io_in_b_37; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_a = io_in_a_38; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_38_io_in_b = io_in_b_38; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_a = io_in_a_39; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_39_io_in_b = io_in_b_39; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_a = io_in_a_40; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_40_io_in_b = io_in_b_40; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_a = io_in_a_41; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_41_io_in_b = io_in_b_41; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_a = io_in_a_42; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_42_io_in_b = io_in_b_42; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_a = io_in_a_43; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_43_io_in_b = io_in_b_43; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_a = io_in_a_44; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_44_io_in_b = io_in_b_44; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_a = io_in_a_45; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_45_io_in_b = io_in_b_45; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_a = io_in_a_46; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_46_io_in_b = io_in_b_46; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_a = io_in_a_47; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_47_io_in_b = io_in_b_47; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_48_clock = clock;
  assign FP_multiplier_10ccs_48_reset = reset;
  assign FP_multiplier_10ccs_48_io_in_a = io_in_a_48; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_48_io_in_b = io_in_b_48; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_49_clock = clock;
  assign FP_multiplier_10ccs_49_reset = reset;
  assign FP_multiplier_10ccs_49_io_in_a = io_in_a_49; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_49_io_in_b = io_in_b_49; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_50_clock = clock;
  assign FP_multiplier_10ccs_50_reset = reset;
  assign FP_multiplier_10ccs_50_io_in_a = io_in_a_50; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_50_io_in_b = io_in_b_50; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_51_clock = clock;
  assign FP_multiplier_10ccs_51_reset = reset;
  assign FP_multiplier_10ccs_51_io_in_a = io_in_a_51; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_51_io_in_b = io_in_b_51; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_52_clock = clock;
  assign FP_multiplier_10ccs_52_reset = reset;
  assign FP_multiplier_10ccs_52_io_in_a = io_in_a_52; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_52_io_in_b = io_in_b_52; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_53_clock = clock;
  assign FP_multiplier_10ccs_53_reset = reset;
  assign FP_multiplier_10ccs_53_io_in_a = io_in_a_53; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_53_io_in_b = io_in_b_53; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_54_clock = clock;
  assign FP_multiplier_10ccs_54_reset = reset;
  assign FP_multiplier_10ccs_54_io_in_a = io_in_a_54; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_54_io_in_b = io_in_b_54; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_55_clock = clock;
  assign FP_multiplier_10ccs_55_reset = reset;
  assign FP_multiplier_10ccs_55_io_in_a = io_in_a_55; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_55_io_in_b = io_in_b_55; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_56_clock = clock;
  assign FP_multiplier_10ccs_56_reset = reset;
  assign FP_multiplier_10ccs_56_io_in_a = io_in_a_56; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_56_io_in_b = io_in_b_56; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_57_clock = clock;
  assign FP_multiplier_10ccs_57_reset = reset;
  assign FP_multiplier_10ccs_57_io_in_a = io_in_a_57; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_57_io_in_b = io_in_b_57; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_58_clock = clock;
  assign FP_multiplier_10ccs_58_reset = reset;
  assign FP_multiplier_10ccs_58_io_in_a = io_in_a_58; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_58_io_in_b = io_in_b_58; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_59_clock = clock;
  assign FP_multiplier_10ccs_59_reset = reset;
  assign FP_multiplier_10ccs_59_io_in_a = io_in_a_59; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_59_io_in_b = io_in_b_59; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_60_clock = clock;
  assign FP_multiplier_10ccs_60_reset = reset;
  assign FP_multiplier_10ccs_60_io_in_a = io_in_a_60; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_60_io_in_b = io_in_b_60; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_61_clock = clock;
  assign FP_multiplier_10ccs_61_reset = reset;
  assign FP_multiplier_10ccs_61_io_in_a = io_in_a_61; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_61_io_in_b = io_in_b_61; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_62_clock = clock;
  assign FP_multiplier_10ccs_62_reset = reset;
  assign FP_multiplier_10ccs_62_io_in_a = io_in_a_62; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_62_io_in_b = io_in_b_62; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_multiplier_10ccs_63_clock = clock;
  assign FP_multiplier_10ccs_63_reset = reset;
  assign FP_multiplier_10ccs_63_io_in_a = io_in_a_63; // @[FloatingPointDesigns.scala 2413:47]
  assign FP_multiplier_10ccs_63_io_in_b = io_in_b_63; // @[FloatingPointDesigns.scala 2414:47]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_1_clock = clock;
  assign FP_adder_13ccs_1_reset = reset;
  assign FP_adder_13ccs_1_io_in_a = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_1_io_in_b = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_2_clock = clock;
  assign FP_adder_13ccs_2_reset = reset;
  assign FP_adder_13ccs_2_io_in_a = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_2_io_in_b = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_3_clock = clock;
  assign FP_adder_13ccs_3_reset = reset;
  assign FP_adder_13ccs_3_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_3_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_4_clock = clock;
  assign FP_adder_13ccs_4_reset = reset;
  assign FP_adder_13ccs_4_io_in_a = FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_4_io_in_b = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_5_clock = clock;
  assign FP_adder_13ccs_5_reset = reset;
  assign FP_adder_13ccs_5_io_in_a = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_5_io_in_b = FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_6_clock = clock;
  assign FP_adder_13ccs_6_reset = reset;
  assign FP_adder_13ccs_6_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_6_io_in_b = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_7_clock = clock;
  assign FP_adder_13ccs_7_reset = reset;
  assign FP_adder_13ccs_7_io_in_a = FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_7_io_in_b = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_8_clock = clock;
  assign FP_adder_13ccs_8_reset = reset;
  assign FP_adder_13ccs_8_io_in_a = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_8_io_in_b = FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_9_clock = clock;
  assign FP_adder_13ccs_9_reset = reset;
  assign FP_adder_13ccs_9_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_9_io_in_b = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_10_clock = clock;
  assign FP_adder_13ccs_10_reset = reset;
  assign FP_adder_13ccs_10_io_in_a = FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_10_io_in_b = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_11_clock = clock;
  assign FP_adder_13ccs_11_reset = reset;
  assign FP_adder_13ccs_11_io_in_a = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_11_io_in_b = FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_12_clock = clock;
  assign FP_adder_13ccs_12_reset = reset;
  assign FP_adder_13ccs_12_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_12_io_in_b = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_13_clock = clock;
  assign FP_adder_13ccs_13_reset = reset;
  assign FP_adder_13ccs_13_io_in_a = FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_13_io_in_b = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_14_clock = clock;
  assign FP_adder_13ccs_14_reset = reset;
  assign FP_adder_13ccs_14_io_in_a = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_14_io_in_b = FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_15_clock = clock;
  assign FP_adder_13ccs_15_reset = reset;
  assign FP_adder_13ccs_15_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_15_io_in_b = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_16_clock = clock;
  assign FP_adder_13ccs_16_reset = reset;
  assign FP_adder_13ccs_16_io_in_a = FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_16_io_in_b = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_17_clock = clock;
  assign FP_adder_13ccs_17_reset = reset;
  assign FP_adder_13ccs_17_io_in_a = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_17_io_in_b = FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_18_clock = clock;
  assign FP_adder_13ccs_18_reset = reset;
  assign FP_adder_13ccs_18_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_18_io_in_b = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_19_clock = clock;
  assign FP_adder_13ccs_19_reset = reset;
  assign FP_adder_13ccs_19_io_in_a = FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_19_io_in_b = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_20_clock = clock;
  assign FP_adder_13ccs_20_reset = reset;
  assign FP_adder_13ccs_20_io_in_a = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_20_io_in_b = FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_21_clock = clock;
  assign FP_adder_13ccs_21_reset = reset;
  assign FP_adder_13ccs_21_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_21_io_in_b = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_22_clock = clock;
  assign FP_adder_13ccs_22_reset = reset;
  assign FP_adder_13ccs_22_io_in_a = FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_22_io_in_b = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_23_clock = clock;
  assign FP_adder_13ccs_23_reset = reset;
  assign FP_adder_13ccs_23_io_in_a = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_23_io_in_b = FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_24_clock = clock;
  assign FP_adder_13ccs_24_reset = reset;
  assign FP_adder_13ccs_24_io_in_a = FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_24_io_in_b = FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_25_clock = clock;
  assign FP_adder_13ccs_25_reset = reset;
  assign FP_adder_13ccs_25_io_in_a = FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_25_io_in_b = FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_26_clock = clock;
  assign FP_adder_13ccs_26_reset = reset;
  assign FP_adder_13ccs_26_io_in_a = FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_26_io_in_b = FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_27_clock = clock;
  assign FP_adder_13ccs_27_reset = reset;
  assign FP_adder_13ccs_27_io_in_a = FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_27_io_in_b = FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_28_clock = clock;
  assign FP_adder_13ccs_28_reset = reset;
  assign FP_adder_13ccs_28_io_in_a = FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_28_io_in_b = FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_29_clock = clock;
  assign FP_adder_13ccs_29_reset = reset;
  assign FP_adder_13ccs_29_io_in_a = FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_29_io_in_b = FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_30_clock = clock;
  assign FP_adder_13ccs_30_reset = reset;
  assign FP_adder_13ccs_30_io_in_a = FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_30_io_in_b = FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_31_clock = clock;
  assign FP_adder_13ccs_31_reset = reset;
  assign FP_adder_13ccs_31_io_in_a = FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_31_io_in_b = FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_32_clock = clock;
  assign FP_adder_13ccs_32_reset = reset;
  assign FP_adder_13ccs_32_io_in_a = FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_32_io_in_b = FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_33_clock = clock;
  assign FP_adder_13ccs_33_reset = reset;
  assign FP_adder_13ccs_33_io_in_a = FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_33_io_in_b = FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_34_clock = clock;
  assign FP_adder_13ccs_34_reset = reset;
  assign FP_adder_13ccs_34_io_in_a = FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_34_io_in_b = FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_35_clock = clock;
  assign FP_adder_13ccs_35_reset = reset;
  assign FP_adder_13ccs_35_io_in_a = FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_35_io_in_b = FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_36_clock = clock;
  assign FP_adder_13ccs_36_reset = reset;
  assign FP_adder_13ccs_36_io_in_a = FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_36_io_in_b = FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_37_clock = clock;
  assign FP_adder_13ccs_37_reset = reset;
  assign FP_adder_13ccs_37_io_in_a = FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_37_io_in_b = FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_38_clock = clock;
  assign FP_adder_13ccs_38_reset = reset;
  assign FP_adder_13ccs_38_io_in_a = FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_38_io_in_b = FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_39_clock = clock;
  assign FP_adder_13ccs_39_reset = reset;
  assign FP_adder_13ccs_39_io_in_a = FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_39_io_in_b = FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_40_clock = clock;
  assign FP_adder_13ccs_40_reset = reset;
  assign FP_adder_13ccs_40_io_in_a = FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_40_io_in_b = FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_41_clock = clock;
  assign FP_adder_13ccs_41_reset = reset;
  assign FP_adder_13ccs_41_io_in_a = FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_41_io_in_b = FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_42_clock = clock;
  assign FP_adder_13ccs_42_reset = reset;
  assign FP_adder_13ccs_42_io_in_a = FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_42_io_in_b = FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_43_clock = clock;
  assign FP_adder_13ccs_43_reset = reset;
  assign FP_adder_13ccs_43_io_in_a = FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_43_io_in_b = FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_44_clock = clock;
  assign FP_adder_13ccs_44_reset = reset;
  assign FP_adder_13ccs_44_io_in_a = FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_44_io_in_b = FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_45_clock = clock;
  assign FP_adder_13ccs_45_reset = reset;
  assign FP_adder_13ccs_45_io_in_a = FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_45_io_in_b = FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_46_clock = clock;
  assign FP_adder_13ccs_46_reset = reset;
  assign FP_adder_13ccs_46_io_in_a = FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_46_io_in_b = FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_47_clock = clock;
  assign FP_adder_13ccs_47_reset = reset;
  assign FP_adder_13ccs_47_io_in_a = FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_47_io_in_b = FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_48_clock = clock;
  assign FP_adder_13ccs_48_reset = reset;
  assign FP_adder_13ccs_48_io_in_a = FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_48_io_in_b = FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_49_clock = clock;
  assign FP_adder_13ccs_49_reset = reset;
  assign FP_adder_13ccs_49_io_in_a = FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_49_io_in_b = FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_50_clock = clock;
  assign FP_adder_13ccs_50_reset = reset;
  assign FP_adder_13ccs_50_io_in_a = FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_50_io_in_b = FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_51_clock = clock;
  assign FP_adder_13ccs_51_reset = reset;
  assign FP_adder_13ccs_51_io_in_a = FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_51_io_in_b = FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_52_clock = clock;
  assign FP_adder_13ccs_52_reset = reset;
  assign FP_adder_13ccs_52_io_in_a = FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_52_io_in_b = FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_53_clock = clock;
  assign FP_adder_13ccs_53_reset = reset;
  assign FP_adder_13ccs_53_io_in_a = FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_53_io_in_b = FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_54_clock = clock;
  assign FP_adder_13ccs_54_reset = reset;
  assign FP_adder_13ccs_54_io_in_a = FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_54_io_in_b = FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_55_clock = clock;
  assign FP_adder_13ccs_55_reset = reset;
  assign FP_adder_13ccs_55_io_in_a = FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_55_io_in_b = FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_56_clock = clock;
  assign FP_adder_13ccs_56_reset = reset;
  assign FP_adder_13ccs_56_io_in_a = FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_56_io_in_b = FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_57_clock = clock;
  assign FP_adder_13ccs_57_reset = reset;
  assign FP_adder_13ccs_57_io_in_a = FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_57_io_in_b = FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_58_clock = clock;
  assign FP_adder_13ccs_58_reset = reset;
  assign FP_adder_13ccs_58_io_in_a = FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_58_io_in_b = FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_59_clock = clock;
  assign FP_adder_13ccs_59_reset = reset;
  assign FP_adder_13ccs_59_io_in_a = FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_59_io_in_b = FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_60_clock = clock;
  assign FP_adder_13ccs_60_reset = reset;
  assign FP_adder_13ccs_60_io_in_a = FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_60_io_in_b = FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_61_clock = clock;
  assign FP_adder_13ccs_61_reset = reset;
  assign FP_adder_13ccs_61_io_in_a = FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_61_io_in_b = FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  assign FP_adder_13ccs_62_clock = clock;
  assign FP_adder_13ccs_62_reset = reset;
  assign FP_adder_13ccs_62_io_in_a = FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2450:43]
  assign FP_adder_13ccs_62_io_in_b = FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2451:43]
  always @(posedge clock) begin
    io_out_s_REG <= FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2468:26]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_s_REG = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FP_subtractor_13ccs(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_clock; // @[FloatingPointDesigns.scala 1650:26]
  wire  FP_adder_reset; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_in_a; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_in_b; // @[FloatingPointDesigns.scala 1650:26]
  wire [31:0] FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1650:26]
  wire  _adjusted_in_b_T_1 = ~io_in_b[31]; // @[FloatingPointDesigns.scala 1653:23]
  FP_adder_13ccs FP_adder ( // @[FloatingPointDesigns.scala 1650:26]
    .clock(FP_adder_clock),
    .reset(FP_adder_reset),
    .io_in_a(FP_adder_io_in_a),
    .io_in_b(FP_adder_io_in_b),
    .io_out_s(FP_adder_io_out_s)
  );
  assign io_out_s = FP_adder_io_out_s; // @[FloatingPointDesigns.scala 1657:14]
  assign FP_adder_clock = clock;
  assign FP_adder_reset = reset;
  assign FP_adder_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 1655:22]
  assign FP_adder_io_in_b = {_adjusted_in_b_T_1,io_in_b[30:0]}; // @[FloatingPointDesigns.scala 1653:41]
endmodule
module FP_square_root_newfpu(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 1878:65]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 1878:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 1879:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 1879:50]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 1879:50]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1879:50]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 1879:50]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 1879:50]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1879:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 1947:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 1947:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 1947:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 1947:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 1947:29]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 1862:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 1859:46 1860:14 1862:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1856:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 1869:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_4; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_5; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_6; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_8; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_9; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] x_n_10; // @[FloatingPointDesigns.scala 1871:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_4; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_5; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_6; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_7; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_8; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_9; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_10; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] a_2_11; // @[FloatingPointDesigns.scala 1872:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_1_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_0_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_0; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_1; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_2; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_3; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_4; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_5; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_6; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_7; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage1_regs_2_1_8; // @[FloatingPointDesigns.scala 1873:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_0_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_1_1_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_0_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_0; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_1; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_2; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_3; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_4; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_5; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_6; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_7; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage2_regs_2_1_8; // @[FloatingPointDesigns.scala 1874:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_0_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_1_1_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_0_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_0; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_1; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_2; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_3; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_4; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_5; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_6; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_7; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_8; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_9; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_10; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage3_regs_2_1_11; // @[FloatingPointDesigns.scala 1875:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_0; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_1; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_2; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_3; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_4; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_5; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_6; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_7; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_1_1_8; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_0; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_1; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_2; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_3; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_4; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_5; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_6; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_7; // @[FloatingPointDesigns.scala 1876:30]
  reg [31:0] stage4_regs_2_1_8; // @[FloatingPointDesigns.scala 1876:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 1901:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 1901:82]
  wire [31:0] _GEN_139 = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1871:22 1908:28 1909:26]
  wire [31:0] _GEN_215 = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 1871:22 1908:28 1909:26]
  wire [7:0] _restore_a_T_3 = stage4_regs_2_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 1946:106]
  wire [8:0] _restore_a_T_4 = {stage4_regs_2_1_8[31],_restore_a_T_3}; // @[FloatingPointDesigns.scala 1946:55]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 1878:65]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 1879:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 1879:50]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 1879:50]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 1947:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  assign io_out_s = {{1'd0}, multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1951:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 1905:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 1906:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 1918:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 1919:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 1936:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 1937:34]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1914:48]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1915:48]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 1918:34]
  assign FP_multiplier_10ccs_4_io_in_b = {1'h0,stage1_regs_1_1_8[30:0]}; // @[FloatingPointDesigns.scala 1919:46]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,stage3_regs_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 1936:46]
  assign FP_multiplier_10ccs_5_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1937:34]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1914:48]
  assign FP_multiplier_10ccs_6_io_in_b = {1'h0,FP_multiplier_10ccs_5_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1915:48]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 1918:34]
  assign FP_multiplier_10ccs_7_io_in_b = {1'h0,stage1_regs_2_1_8[30:0]}; // @[FloatingPointDesigns.scala 1919:46]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = {1'h0,stage3_regs_2_0_11[30:0]}; // @[FloatingPointDesigns.scala 1936:46]
  assign FP_multiplier_10ccs_8_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 1937:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1857:26 1858:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 1928:31]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1857:26 1858:16]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 1928:31]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1857:26 1858:16]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 1928:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_8_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 1949:37]
  assign multiplier4_io_in_b = {_restore_a_T_4,stage4_regs_2_1_8[22:0]}; // @[FloatingPointDesigns.scala 1946:113]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_0 <= result;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_1 <= stage1_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_2 <= stage2_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_4 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_4 <= _GEN_139;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_5 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_5 <= stage1_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_6 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_6 <= stage2_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_8 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_8 <= _GEN_215;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_9 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_9 <= stage1_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1871:22]
      x_n_10 <= 32'h0; // @[FloatingPointDesigns.scala 1871:22]
    end else begin
      x_n_10 <= stage2_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_0 <= _a_2_0_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_1 <= stage1_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_2 <= stage2_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_3 <= stage3_regs_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_4 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_4 <= stage4_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_5 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_5 <= stage1_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_6 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_6 <= stage2_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_7 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_7 <= stage3_regs_1_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_8 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_8 <= stage4_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_9 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_9 <= stage1_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_10 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_10 <= stage2_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1872:22]
      a_2_11 <= 32'h0; // @[FloatingPointDesigns.scala 1872:22]
    end else begin
      a_2_11 <= stage3_regs_2_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_0 <= x_n_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_1 <= stage1_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_2 <= stage1_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_3 <= stage1_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_4 <= stage1_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_5 <= stage1_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_6 <= stage1_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_7 <= stage1_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_0_8 <= stage1_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_0 <= a_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_1 <= stage1_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_2 <= stage1_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_3 <= stage1_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_4 <= stage1_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_5 <= stage1_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_6 <= stage1_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_7 <= stage1_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_0_1_8 <= stage1_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_0 <= x_n_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_1 <= stage1_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_2 <= stage1_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_3 <= stage1_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_4 <= stage1_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_5 <= stage1_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_6 <= stage1_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_7 <= stage1_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_0_8 <= stage1_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_0 <= a_2_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_1 <= stage1_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_2 <= stage1_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_3 <= stage1_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_4 <= stage1_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_5 <= stage1_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_6 <= stage1_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_7 <= stage1_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_1_1_8 <= stage1_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_0 <= x_n_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_1 <= stage1_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_2 <= stage1_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_3 <= stage1_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_4 <= stage1_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_5 <= stage1_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_6 <= stage1_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_7 <= stage1_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_0_8 <= stage1_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_0 <= a_2_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_1 <= stage1_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_2 <= stage1_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_3 <= stage1_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_4 <= stage1_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_5 <= stage1_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_6 <= stage1_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_7 <= stage1_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1873:30]
      stage1_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1873:30]
    end else begin
      stage1_regs_2_1_8 <= stage1_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_0 <= x_n_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_1 <= stage2_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_2 <= stage2_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_3 <= stage2_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_4 <= stage2_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_5 <= stage2_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_6 <= stage2_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_7 <= stage2_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_0_8 <= stage2_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_0 <= a_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_1 <= stage2_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_2 <= stage2_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_3 <= stage2_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_4 <= stage2_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_5 <= stage2_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_6 <= stage2_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_7 <= stage2_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_0_1_8 <= stage2_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_0 <= x_n_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_1 <= stage2_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_2 <= stage2_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_3 <= stage2_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_4 <= stage2_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_5 <= stage2_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_6 <= stage2_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_7 <= stage2_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_0_8 <= stage2_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_0 <= a_2_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_1 <= stage2_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_2 <= stage2_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_3 <= stage2_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_4 <= stage2_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_5 <= stage2_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_6 <= stage2_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_7 <= stage2_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_1_1_8 <= stage2_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_0 <= x_n_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_1 <= stage2_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_2 <= stage2_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_3 <= stage2_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_4 <= stage2_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_5 <= stage2_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_6 <= stage2_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_7 <= stage2_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_0_8 <= stage2_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_0 <= a_2_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_1 <= stage2_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_2 <= stage2_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_3 <= stage2_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_4 <= stage2_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_5 <= stage2_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_6 <= stage2_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_7 <= stage2_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1874:30]
      stage2_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1874:30]
    end else begin
      stage2_regs_2_1_8 <= stage2_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_0 <= x_n_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_1 <= stage3_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_2 <= stage3_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_3 <= stage3_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_4 <= stage3_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_5 <= stage3_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_6 <= stage3_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_7 <= stage3_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_8 <= stage3_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_9 <= stage3_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_10 <= stage3_regs_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_0_11 <= stage3_regs_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_0 <= a_2_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_1 <= stage3_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_2 <= stage3_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_3 <= stage3_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_4 <= stage3_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_5 <= stage3_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_6 <= stage3_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_7 <= stage3_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_8 <= stage3_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_9 <= stage3_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_10 <= stage3_regs_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_0_1_11 <= stage3_regs_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_0 <= x_n_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_1 <= stage3_regs_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_2 <= stage3_regs_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_3 <= stage3_regs_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_4 <= stage3_regs_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_5 <= stage3_regs_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_6 <= stage3_regs_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_7 <= stage3_regs_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_8 <= stage3_regs_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_9 <= stage3_regs_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_10 <= stage3_regs_1_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_0_11 <= stage3_regs_1_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_0 <= a_2_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_1 <= stage3_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_2 <= stage3_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_3 <= stage3_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_4 <= stage3_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_5 <= stage3_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_6 <= stage3_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_7 <= stage3_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_8 <= stage3_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_9 <= stage3_regs_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_10 <= stage3_regs_1_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_1_1_11 <= stage3_regs_1_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_0 <= x_n_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_1 <= stage3_regs_2_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_2 <= stage3_regs_2_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_3 <= stage3_regs_2_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_4 <= stage3_regs_2_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_5 <= stage3_regs_2_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_6 <= stage3_regs_2_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_7 <= stage3_regs_2_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_8 <= stage3_regs_2_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_9 <= stage3_regs_2_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_10 <= stage3_regs_2_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_0_11 <= stage3_regs_2_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_0 <= a_2_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_1 <= stage3_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_2 <= stage3_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_3 <= stage3_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_4 <= stage3_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_5 <= stage3_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_6 <= stage3_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_7 <= stage3_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_8 <= stage3_regs_2_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_9 <= stage3_regs_2_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_10 <= stage3_regs_2_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1875:30]
      stage3_regs_2_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 1875:30]
    end else begin
      stage3_regs_2_1_11 <= stage3_regs_2_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_0 <= a_2_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_1 <= stage4_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_2 <= stage4_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_3 <= stage4_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_4 <= stage4_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_5 <= stage4_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_6 <= stage4_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_7 <= stage4_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_0_1_8 <= stage4_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_0 <= a_2_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_1 <= stage4_regs_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_2 <= stage4_regs_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_3 <= stage4_regs_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_4 <= stage4_regs_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_5 <= stage4_regs_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_6 <= stage4_regs_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_7 <= stage4_regs_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_1_1_8 <= stage4_regs_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_0 <= a_2_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_1 <= stage4_regs_2_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_2 <= stage4_regs_2_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_3 <= stage4_regs_2_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_4 <= stage4_regs_2_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_5 <= stage4_regs_2_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_6 <= stage4_regs_2_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_7 <= stage4_regs_2_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 1876:30]
      stage4_regs_2_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 1876:30]
    end else begin
      stage4_regs_2_1_8 <= stage4_regs_2_1_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  x_n_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  x_n_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  x_n_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  x_n_8 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  x_n_9 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  x_n_10 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  a_2_0 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  a_2_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  a_2_2 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  a_2_3 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  a_2_4 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  a_2_5 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  a_2_6 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  a_2_7 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  a_2_8 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  a_2_9 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  a_2_10 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  a_2_11 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  stage1_regs_1_0_0 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  stage1_regs_1_0_1 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  stage1_regs_1_0_2 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  stage1_regs_1_0_3 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  stage1_regs_1_0_4 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  stage1_regs_1_0_5 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  stage1_regs_1_0_6 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  stage1_regs_1_0_7 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  stage1_regs_1_0_8 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  stage1_regs_1_1_0 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  stage1_regs_1_1_1 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  stage1_regs_1_1_2 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  stage1_regs_1_1_3 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  stage1_regs_1_1_4 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  stage1_regs_1_1_5 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  stage1_regs_1_1_6 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  stage1_regs_1_1_7 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  stage1_regs_1_1_8 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  stage1_regs_2_0_0 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  stage1_regs_2_0_1 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  stage1_regs_2_0_2 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  stage1_regs_2_0_3 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  stage1_regs_2_0_4 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  stage1_regs_2_0_5 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  stage1_regs_2_0_6 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  stage1_regs_2_0_7 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  stage1_regs_2_0_8 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  stage1_regs_2_1_0 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  stage1_regs_2_1_1 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  stage1_regs_2_1_2 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  stage1_regs_2_1_3 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  stage1_regs_2_1_4 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  stage1_regs_2_1_5 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  stage1_regs_2_1_6 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  stage1_regs_2_1_7 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  stage1_regs_2_1_8 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  stage2_regs_1_0_0 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  stage2_regs_1_0_1 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  stage2_regs_1_0_2 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  stage2_regs_1_0_3 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  stage2_regs_1_0_4 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  stage2_regs_1_0_5 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  stage2_regs_1_0_6 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  stage2_regs_1_0_7 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  stage2_regs_1_0_8 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  stage2_regs_1_1_0 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  stage2_regs_1_1_1 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  stage2_regs_1_1_2 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  stage2_regs_1_1_3 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  stage2_regs_1_1_4 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  stage2_regs_1_1_5 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  stage2_regs_1_1_6 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  stage2_regs_1_1_7 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  stage2_regs_1_1_8 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  stage2_regs_2_0_0 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage2_regs_2_0_1 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage2_regs_2_0_2 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage2_regs_2_0_3 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage2_regs_2_0_4 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage2_regs_2_0_5 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage2_regs_2_0_6 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage2_regs_2_0_7 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage2_regs_2_0_8 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage2_regs_2_1_0 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage2_regs_2_1_1 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage2_regs_2_1_2 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage2_regs_2_1_3 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage2_regs_2_1_4 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage2_regs_2_1_5 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage2_regs_2_1_6 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage2_regs_2_1_7 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage2_regs_2_1_8 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage3_regs_1_0_0 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage3_regs_1_0_1 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage3_regs_1_0_2 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage3_regs_1_0_3 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage3_regs_1_0_4 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage3_regs_1_0_5 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage3_regs_1_0_6 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage3_regs_1_0_7 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage3_regs_1_0_8 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage3_regs_1_0_9 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage3_regs_1_0_10 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage3_regs_1_0_11 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage3_regs_1_1_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage3_regs_1_1_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage3_regs_1_1_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage3_regs_1_1_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage3_regs_1_1_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage3_regs_1_1_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage3_regs_1_1_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage3_regs_1_1_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage3_regs_1_1_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage3_regs_1_1_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage3_regs_1_1_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage3_regs_1_1_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage3_regs_2_0_0 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage3_regs_2_0_1 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage3_regs_2_0_2 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage3_regs_2_0_3 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage3_regs_2_0_4 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage3_regs_2_0_5 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage3_regs_2_0_6 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage3_regs_2_0_7 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage3_regs_2_0_8 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage3_regs_2_0_9 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage3_regs_2_0_10 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage3_regs_2_0_11 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage3_regs_2_1_0 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage3_regs_2_1_1 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage3_regs_2_1_2 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage3_regs_2_1_3 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage3_regs_2_1_4 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage3_regs_2_1_5 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage3_regs_2_1_6 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage3_regs_2_1_7 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage3_regs_2_1_8 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  stage3_regs_2_1_9 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  stage3_regs_2_1_10 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  stage3_regs_2_1_11 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  stage4_regs_1_1_0 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  stage4_regs_1_1_1 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  stage4_regs_1_1_2 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  stage4_regs_1_1_3 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  stage4_regs_1_1_4 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  stage4_regs_1_1_5 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  stage4_regs_1_1_6 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  stage4_regs_1_1_7 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  stage4_regs_1_1_8 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  stage4_regs_2_1_0 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  stage4_regs_2_1_1 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  stage4_regs_2_1_2 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  stage4_regs_2_1_3 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  stage4_regs_2_1_4 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  stage4_regs_2_1_5 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  stage4_regs_2_1_6 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  stage4_regs_2_1_7 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  stage4_regs_2_1_8 = _RAND_227[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hqr5(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b,
  output [31:0] io_out_s
);
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2512:23]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2512:23]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2512:23]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2512:23]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2512:23]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 2513:28]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 2513:28]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2513:28]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2513:28]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2513:28]
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2512:23]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 2513:28]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  assign io_out_s = io_in_a[31] ? FP_subtractor_13ccs_io_out_s : FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2521:24 2522:14 2524:14]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2515:16]
  assign FP_adder_13ccs_io_in_b = io_in_b; // @[FloatingPointDesigns.scala 2516:16]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2518:21]
  assign FP_subtractor_13ccs_io_in_b = io_in_b; // @[FloatingPointDesigns.scala 2519:21]
endmodule
module FP_reciprocal_newfpu(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
`endif // RANDOMIZE_REG_INIT
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2007:65]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2007:65]
  wire  FP_subtractor_13ccs_clock; // @[FloatingPointDesigns.scala 2008:50]
  wire  FP_subtractor_13ccs_reset; // @[FloatingPointDesigns.scala 2008:50]
  wire [31:0] FP_subtractor_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2008:50]
  wire [31:0] FP_subtractor_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2008:50]
  wire [31:0] FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2008:50]
  wire  multiplier4_clock; // @[FloatingPointDesigns.scala 2087:29]
  wire  multiplier4_reset; // @[FloatingPointDesigns.scala 2087:29]
  wire [31:0] multiplier4_io_in_a; // @[FloatingPointDesigns.scala 2087:29]
  wire [31:0] multiplier4_io_in_b; // @[FloatingPointDesigns.scala 2087:29]
  wire [31:0] multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2087:29]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2099:69]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2099:69]
  wire  FP_subtractor_13ccs_1_clock; // @[FloatingPointDesigns.scala 2100:54]
  wire  FP_subtractor_13ccs_1_reset; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2100:54]
  wire  FP_subtractor_13ccs_2_clock; // @[FloatingPointDesigns.scala 2100:54]
  wire  FP_subtractor_13ccs_2_reset; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2100:54]
  wire [31:0] FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2100:54]
  wire [30:0] _number_T_1 = {{1'd0}, io_in_a[30:1]}; // @[FloatingPointDesigns.scala 1992:36]
  wire [30:0] _GEN_0 = io_in_a[30:0] > 31'h7ef477d4 ? 31'h3f7a3bea : _number_T_1; // @[FloatingPointDesigns.scala 1989:46 1990:14 1992:14]
  wire [31:0] number = {{1'd0}, _GEN_0}; // @[FloatingPointDesigns.scala 1984:22]
  wire [31:0] result = 32'h5f3759df - number; // @[FloatingPointDesigns.scala 1999:25]
  reg [31:0] x_n_0; // @[FloatingPointDesigns.scala 2001:22]
  reg [31:0] x_n_1; // @[FloatingPointDesigns.scala 2001:22]
  reg [31:0] x_n_2; // @[FloatingPointDesigns.scala 2001:22]
  reg [31:0] a_2_0; // @[FloatingPointDesigns.scala 2002:22]
  reg [31:0] a_2_1; // @[FloatingPointDesigns.scala 2002:22]
  reg [31:0] a_2_2; // @[FloatingPointDesigns.scala 2002:22]
  reg [31:0] a_2_3; // @[FloatingPointDesigns.scala 2002:22]
  reg [31:0] stage1_regs_0_0_0; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_1; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_2; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_3; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_4; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_5; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_6; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_7; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_0_8; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_0; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_1; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_2; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_3; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_4; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_5; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_6; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_7; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage1_regs_0_1_8; // @[FloatingPointDesigns.scala 2003:30]
  reg [31:0] stage2_regs_0_0_0; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_1; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_2; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_3; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_4; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_5; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_6; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_7; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_0_8; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_0; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_1; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_2; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_3; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_4; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_5; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_6; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_7; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage2_regs_0_1_8; // @[FloatingPointDesigns.scala 2004:30]
  reg [31:0] stage3_regs_0_0_0; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_1; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_2; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_3; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_4; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_5; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_6; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_7; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_8; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_9; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_10; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_0_11; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_0; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_1; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_2; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_3; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_4; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_5; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_6; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_7; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_8; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_9; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_10; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage3_regs_0_1_11; // @[FloatingPointDesigns.scala 2005:30]
  reg [31:0] stage4_regs_0_1_0; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_1; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_2; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_3; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_4; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_5; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_6; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_7; // @[FloatingPointDesigns.scala 2006:30]
  reg [31:0] stage4_regs_0_1_8; // @[FloatingPointDesigns.scala 2006:30]
  wire [7:0] _a_2_0_T_3 = io_in_a[30:23] - 8'h1; // @[FloatingPointDesigns.scala 2032:75]
  wire [31:0] _a_2_0_T_6 = {io_in_a[31],_a_2_0_T_3,io_in_a[22:0]}; // @[FloatingPointDesigns.scala 2032:82]
  reg [31:0] a_2_isr_to_r; // @[FloatingPointDesigns.scala 2077:31]
  reg [31:0] transition_regs_0; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_1; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_2; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_3; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_4; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_5; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_6; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_7; // @[FloatingPointDesigns.scala 2078:34]
  reg [31:0] transition_regs_8; // @[FloatingPointDesigns.scala 2078:34]
  wire [7:0] _a_2_isr_to_r_T_3 = stage4_regs_0_1_8[30:23] + 8'h1; // @[FloatingPointDesigns.scala 2080:115]
  wire [31:0] _a_2_isr_to_r_T_6 = {stage4_regs_0_1_8[31],_a_2_isr_to_r_T_3,stage4_regs_0_1_8[22:0]}; // @[FloatingPointDesigns.scala 2080:122]
  reg [31:0] x_n_r_0; // @[FloatingPointDesigns.scala 2094:24]
  reg [31:0] x_n_r_1; // @[FloatingPointDesigns.scala 2094:24]
  reg [31:0] x_n_r_3; // @[FloatingPointDesigns.scala 2094:24]
  reg [31:0] x_n_r_4; // @[FloatingPointDesigns.scala 2094:24]
  reg [31:0] a_2_r_0; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] a_2_r_1; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] a_2_r_2; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] a_2_r_3; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] a_2_r_4; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] a_2_r_5; // @[FloatingPointDesigns.scala 2095:24]
  reg [31:0] stage1_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage1_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2096:32]
  reg [31:0] stage2_regs_r_0_0_0; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_1; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_2; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_3; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_4; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_5; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_6; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_7; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_8; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_9; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_10; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_0_11; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_9; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_10; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_0_1_11; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_0; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_1; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_2; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_3; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_4; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_5; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_6; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_7; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_8; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_9; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_10; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_0_11; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_9; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_10; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage2_regs_r_1_1_11; // @[FloatingPointDesigns.scala 2097:32]
  reg [31:0] stage3_regs_r_0_1_0; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_1; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_2; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_3; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_4; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_5; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_6; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_7; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_0_1_8; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_0; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_1; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_2; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_3; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_4; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_5; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_6; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_7; // @[FloatingPointDesigns.scala 2098:32]
  reg [31:0] stage3_regs_r_1_1_8; // @[FloatingPointDesigns.scala 2098:32]
  wire [31:0] _GEN_133 = multiplier4_io_out_s; // @[FloatingPointDesigns.scala 2094:24 2119:28 2120:28]
  wire [31:0] _GEN_189 = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2094:24 2128:28 2129:28]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2007:65]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2007:65]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2007:65]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs ( // @[FloatingPointDesigns.scala 2008:50]
    .clock(FP_subtractor_13ccs_clock),
    .reset(FP_subtractor_13ccs_reset),
    .io_in_a(FP_subtractor_13ccs_io_in_a),
    .io_in_b(FP_subtractor_13ccs_io_in_b),
    .io_out_s(FP_subtractor_13ccs_io_out_s)
  );
  FP_multiplier_10ccs multiplier4 ( // @[FloatingPointDesigns.scala 2087:29]
    .clock(multiplier4_clock),
    .reset(multiplier4_reset),
    .io_in_a(multiplier4_io_in_a),
    .io_in_b(multiplier4_io_in_b),
    .io_out_s(multiplier4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2099:69]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2099:69]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2099:69]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2099:69]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_1 ( // @[FloatingPointDesigns.scala 2100:54]
    .clock(FP_subtractor_13ccs_1_clock),
    .reset(FP_subtractor_13ccs_1_reset),
    .io_in_a(FP_subtractor_13ccs_1_io_in_a),
    .io_in_b(FP_subtractor_13ccs_1_io_in_b),
    .io_out_s(FP_subtractor_13ccs_1_io_out_s)
  );
  FP_subtractor_13ccs FP_subtractor_13ccs_2 ( // @[FloatingPointDesigns.scala 2100:54]
    .clock(FP_subtractor_13ccs_2_clock),
    .reset(FP_subtractor_13ccs_2_reset),
    .io_in_a(FP_subtractor_13ccs_2_io_in_a),
    .io_in_b(FP_subtractor_13ccs_2_io_in_b),
    .io_out_s(FP_subtractor_13ccs_2_io_out_s)
  );
  assign io_out_s = {stage3_regs_r_1_1_8[31],FP_multiplier_10ccs_6_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2156:58]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2036:48]
  assign FP_multiplier_10ccs_io_in_b = {1'h0,result[30:0]}; // @[FloatingPointDesigns.scala 2037:48]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2049:34]
  assign FP_multiplier_10ccs_1_io_in_b = {1'h0,stage1_regs_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2050:46]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = {1'h0,stage3_regs_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2067:46]
  assign FP_multiplier_10ccs_2_io_in_b = FP_subtractor_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2068:34]
  assign FP_subtractor_13ccs_clock = clock;
  assign FP_subtractor_13ccs_reset = reset;
  assign FP_subtractor_13ccs_io_in_a = 32'h3fc00000; // @[FloatingPointDesigns.scala 1985:26 1986:16]
  assign FP_subtractor_13ccs_io_in_b = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2059:31]
  assign multiplier4_clock = clock;
  assign multiplier4_reset = reset;
  assign multiplier4_io_in_a = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2089:37]
  assign multiplier4_io_in_b = {1'h0,FP_multiplier_10ccs_2_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2090:37]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = {1'h0,multiplier4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2125:50]
  assign FP_multiplier_10ccs_3_io_in_b = {1'h0,transition_regs_8[30:0]}; // @[FloatingPointDesigns.scala 2126:50]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = {1'h0,stage2_regs_r_0_0_11[30:0]}; // @[FloatingPointDesigns.scala 2147:48]
  assign FP_multiplier_10ccs_4_io_in_b = FP_subtractor_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2148:36]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = {1'h0,FP_multiplier_10ccs_4_io_out_s[30:0]}; // @[FloatingPointDesigns.scala 2134:50]
  assign FP_multiplier_10ccs_5_io_in_b = {1'h0,stage3_regs_r_0_1_8[30:0]}; // @[FloatingPointDesigns.scala 2135:50]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = {1'h0,stage2_regs_r_1_0_11[30:0]}; // @[FloatingPointDesigns.scala 2147:48]
  assign FP_multiplier_10ccs_6_io_in_b = FP_subtractor_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2148:36]
  assign FP_subtractor_13ccs_1_clock = clock;
  assign FP_subtractor_13ccs_1_reset = reset;
  assign FP_subtractor_13ccs_1_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 1987:19 1988:9]
  assign FP_subtractor_13ccs_1_io_in_b = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2139:33]
  assign FP_subtractor_13ccs_2_clock = clock;
  assign FP_subtractor_13ccs_2_reset = reset;
  assign FP_subtractor_13ccs_2_io_in_a = 32'h40000000; // @[FloatingPointDesigns.scala 1987:19 1988:9]
  assign FP_subtractor_13ccs_2_io_in_b = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2139:33]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2001:22]
      x_n_0 <= 32'h0; // @[FloatingPointDesigns.scala 2001:22]
    end else begin
      x_n_0 <= result;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:22]
      x_n_1 <= 32'h0; // @[FloatingPointDesigns.scala 2001:22]
    end else begin
      x_n_1 <= stage1_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2001:22]
      x_n_2 <= 32'h0; // @[FloatingPointDesigns.scala 2001:22]
    end else begin
      x_n_2 <= stage2_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:22]
      a_2_0 <= 32'h0; // @[FloatingPointDesigns.scala 2002:22]
    end else begin
      a_2_0 <= _a_2_0_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:22]
      a_2_1 <= 32'h0; // @[FloatingPointDesigns.scala 2002:22]
    end else begin
      a_2_1 <= stage1_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:22]
      a_2_2 <= 32'h0; // @[FloatingPointDesigns.scala 2002:22]
    end else begin
      a_2_2 <= stage2_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2002:22]
      a_2_3 <= 32'h0; // @[FloatingPointDesigns.scala 2002:22]
    end else begin
      a_2_3 <= stage3_regs_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_0 <= x_n_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_1 <= stage1_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_2 <= stage1_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_3 <= stage1_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_4 <= stage1_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_5 <= stage1_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_6 <= stage1_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_7 <= stage1_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_0_8 <= stage1_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_0 <= a_2_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_1 <= stage1_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_2 <= stage1_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_3 <= stage1_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_4 <= stage1_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_5 <= stage1_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_6 <= stage1_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_7 <= stage1_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2003:30]
      stage1_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2003:30]
    end else begin
      stage1_regs_0_1_8 <= stage1_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_0 <= x_n_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_1 <= stage2_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_2 <= stage2_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_3 <= stage2_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_4 <= stage2_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_5 <= stage2_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_6 <= stage2_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_7 <= stage2_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_0_8 <= stage2_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_0 <= a_2_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_1 <= stage2_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_2 <= stage2_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_3 <= stage2_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_4 <= stage2_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_5 <= stage2_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_6 <= stage2_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_7 <= stage2_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2004:30]
      stage2_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2004:30]
    end else begin
      stage2_regs_0_1_8 <= stage2_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_0 <= x_n_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_1 <= stage3_regs_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_2 <= stage3_regs_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_3 <= stage3_regs_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_4 <= stage3_regs_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_5 <= stage3_regs_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_6 <= stage3_regs_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_7 <= stage3_regs_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_8 <= stage3_regs_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_9 <= stage3_regs_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_10 <= stage3_regs_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_0_11 <= stage3_regs_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_0 <= a_2_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_1 <= stage3_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_2 <= stage3_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_3 <= stage3_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_4 <= stage3_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_5 <= stage3_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_6 <= stage3_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_7 <= stage3_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_8 <= stage3_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_9 <= stage3_regs_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_10 <= stage3_regs_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2005:30]
      stage3_regs_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2005:30]
    end else begin
      stage3_regs_0_1_11 <= stage3_regs_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_0 <= a_2_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_1 <= stage4_regs_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_2 <= stage4_regs_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_3 <= stage4_regs_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_4 <= stage4_regs_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_5 <= stage4_regs_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_6 <= stage4_regs_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_7 <= stage4_regs_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2006:30]
      stage4_regs_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2006:30]
    end else begin
      stage4_regs_0_1_8 <= stage4_regs_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2077:31]
      a_2_isr_to_r <= 32'h0; // @[FloatingPointDesigns.scala 2077:31]
    end else begin
      a_2_isr_to_r <= _a_2_isr_to_r_T_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_0 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_0 <= a_2_isr_to_r;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_1 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_1 <= transition_regs_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_2 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_2 <= transition_regs_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_3 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_3 <= transition_regs_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_4 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_4 <= transition_regs_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_5 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_5 <= transition_regs_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_6 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_6 <= transition_regs_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_7 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_7 <= transition_regs_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2078:34]
      transition_regs_8 <= 32'h0; // @[FloatingPointDesigns.scala 2078:34]
    end else begin
      transition_regs_8 <= transition_regs_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:24]
      x_n_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2094:24]
    end else begin
      x_n_r_0 <= _GEN_133;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:24]
      x_n_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2094:24]
    end else begin
      x_n_r_1 <= stage1_regs_r_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:24]
      x_n_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2094:24]
    end else begin
      x_n_r_3 <= _GEN_189;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2094:24]
      x_n_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2094:24]
    end else begin
      x_n_r_4 <= stage1_regs_r_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_0 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_0 <= transition_regs_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_1 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_1 <= stage1_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_2 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_2 <= stage2_regs_r_0_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_3 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_3 <= stage3_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_4 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_4 <= stage1_regs_r_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2095:24]
      a_2_r_5 <= 32'h0; // @[FloatingPointDesigns.scala 2095:24]
    end else begin
      a_2_r_5 <= stage2_regs_r_1_1_11;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_0 <= x_n_r_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_1 <= stage1_regs_r_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_2 <= stage1_regs_r_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_3 <= stage1_regs_r_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_4 <= stage1_regs_r_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_5 <= stage1_regs_r_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_6 <= stage1_regs_r_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_7 <= stage1_regs_r_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_0_8 <= stage1_regs_r_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_0 <= a_2_r_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_1 <= stage1_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_2 <= stage1_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_3 <= stage1_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_4 <= stage1_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_5 <= stage1_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_6 <= stage1_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_7 <= stage1_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_0_1_8 <= stage1_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_0 <= x_n_r_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_1 <= stage1_regs_r_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_2 <= stage1_regs_r_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_3 <= stage1_regs_r_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_4 <= stage1_regs_r_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_5 <= stage1_regs_r_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_6 <= stage1_regs_r_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_7 <= stage1_regs_r_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_0_8 <= stage1_regs_r_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_0 <= a_2_r_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_1 <= stage1_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_2 <= stage1_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_3 <= stage1_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_4 <= stage1_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_5 <= stage1_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_6 <= stage1_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_7 <= stage1_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2096:32]
      stage1_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2096:32]
    end else begin
      stage1_regs_r_1_1_8 <= stage1_regs_r_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_0 <= x_n_r_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_1 <= stage2_regs_r_0_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_2 <= stage2_regs_r_0_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_3 <= stage2_regs_r_0_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_4 <= stage2_regs_r_0_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_5 <= stage2_regs_r_0_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_6 <= stage2_regs_r_0_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_7 <= stage2_regs_r_0_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_8 <= stage2_regs_r_0_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_9 <= stage2_regs_r_0_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_10 <= stage2_regs_r_0_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_0_11 <= stage2_regs_r_0_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_0 <= a_2_r_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_1 <= stage2_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_2 <= stage2_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_3 <= stage2_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_4 <= stage2_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_5 <= stage2_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_6 <= stage2_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_7 <= stage2_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_8 <= stage2_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_9 <= stage2_regs_r_0_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_10 <= stage2_regs_r_0_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_0_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_0_1_11 <= stage2_regs_r_0_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_0 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_0 <= x_n_r_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_1 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_1 <= stage2_regs_r_1_0_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_2 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_2 <= stage2_regs_r_1_0_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_3 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_3 <= stage2_regs_r_1_0_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_4 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_4 <= stage2_regs_r_1_0_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_5 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_5 <= stage2_regs_r_1_0_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_6 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_6 <= stage2_regs_r_1_0_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_7 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_7 <= stage2_regs_r_1_0_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_8 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_8 <= stage2_regs_r_1_0_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_9 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_9 <= stage2_regs_r_1_0_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_10 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_10 <= stage2_regs_r_1_0_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_0_11 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_0_11 <= stage2_regs_r_1_0_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_0 <= a_2_r_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_1 <= stage2_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_2 <= stage2_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_3 <= stage2_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_4 <= stage2_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_5 <= stage2_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_6 <= stage2_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_7 <= stage2_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_8 <= stage2_regs_r_1_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_9 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_9 <= stage2_regs_r_1_1_8;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_10 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_10 <= stage2_regs_r_1_1_9;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2097:32]
      stage2_regs_r_1_1_11 <= 32'h0; // @[FloatingPointDesigns.scala 2097:32]
    end else begin
      stage2_regs_r_1_1_11 <= stage2_regs_r_1_1_10;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_0 <= a_2_r_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_1 <= stage3_regs_r_0_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_2 <= stage3_regs_r_0_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_3 <= stage3_regs_r_0_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_4 <= stage3_regs_r_0_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_5 <= stage3_regs_r_0_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_6 <= stage3_regs_r_0_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_7 <= stage3_regs_r_0_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_0_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_0_1_8 <= stage3_regs_r_0_1_7;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_0 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_0 <= a_2_r_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_1 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_1 <= stage3_regs_r_1_1_0;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_2 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_2 <= stage3_regs_r_1_1_1;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_3 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_3 <= stage3_regs_r_1_1_2;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_4 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_4 <= stage3_regs_r_1_1_3;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_5 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_5 <= stage3_regs_r_1_1_4;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_6 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_6 <= stage3_regs_r_1_1_5;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_7 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_7 <= stage3_regs_r_1_1_6;
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2098:32]
      stage3_regs_r_1_1_8 <= 32'h0; // @[FloatingPointDesigns.scala 2098:32]
    end else begin
      stage3_regs_r_1_1_8 <= stage3_regs_r_1_1_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  x_n_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  x_n_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  x_n_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  a_2_0 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  a_2_1 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  a_2_2 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  a_2_3 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  stage1_regs_0_0_0 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  stage1_regs_0_0_1 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  stage1_regs_0_0_2 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  stage1_regs_0_0_3 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  stage1_regs_0_0_4 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  stage1_regs_0_0_5 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  stage1_regs_0_0_6 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  stage1_regs_0_0_7 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  stage1_regs_0_0_8 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  stage1_regs_0_1_0 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  stage1_regs_0_1_1 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  stage1_regs_0_1_2 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  stage1_regs_0_1_3 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  stage1_regs_0_1_4 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  stage1_regs_0_1_5 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  stage1_regs_0_1_6 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  stage1_regs_0_1_7 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  stage1_regs_0_1_8 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  stage2_regs_0_0_0 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  stage2_regs_0_0_1 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  stage2_regs_0_0_2 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  stage2_regs_0_0_3 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  stage2_regs_0_0_4 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  stage2_regs_0_0_5 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  stage2_regs_0_0_6 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  stage2_regs_0_0_7 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  stage2_regs_0_0_8 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  stage2_regs_0_1_0 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  stage2_regs_0_1_1 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  stage2_regs_0_1_2 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  stage2_regs_0_1_3 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  stage2_regs_0_1_4 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  stage2_regs_0_1_5 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  stage2_regs_0_1_6 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  stage2_regs_0_1_7 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  stage2_regs_0_1_8 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  stage3_regs_0_0_0 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  stage3_regs_0_0_1 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  stage3_regs_0_0_2 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  stage3_regs_0_0_3 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  stage3_regs_0_0_4 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  stage3_regs_0_0_5 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  stage3_regs_0_0_6 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  stage3_regs_0_0_7 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  stage3_regs_0_0_8 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  stage3_regs_0_0_9 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  stage3_regs_0_0_10 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  stage3_regs_0_0_11 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  stage3_regs_0_1_0 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  stage3_regs_0_1_1 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  stage3_regs_0_1_2 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  stage3_regs_0_1_3 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  stage3_regs_0_1_4 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  stage3_regs_0_1_5 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  stage3_regs_0_1_6 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  stage3_regs_0_1_7 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  stage3_regs_0_1_8 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  stage3_regs_0_1_9 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  stage3_regs_0_1_10 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  stage3_regs_0_1_11 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  stage4_regs_0_1_0 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  stage4_regs_0_1_1 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  stage4_regs_0_1_2 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  stage4_regs_0_1_3 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  stage4_regs_0_1_4 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  stage4_regs_0_1_5 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  stage4_regs_0_1_6 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  stage4_regs_0_1_7 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  stage4_regs_0_1_8 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  a_2_isr_to_r = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  transition_regs_0 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  transition_regs_1 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  transition_regs_2 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  transition_regs_3 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  transition_regs_4 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  transition_regs_5 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  transition_regs_6 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  transition_regs_7 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  transition_regs_8 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  x_n_r_0 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  x_n_r_1 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  x_n_r_3 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  x_n_r_4 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  a_2_r_0 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  a_2_r_1 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  a_2_r_2 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  a_2_r_3 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  a_2_r_4 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  a_2_r_5 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  stage1_regs_r_0_0_0 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  stage1_regs_r_0_0_1 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  stage1_regs_r_0_0_2 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  stage1_regs_r_0_0_3 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  stage1_regs_r_0_0_4 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  stage1_regs_r_0_0_5 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  stage1_regs_r_0_0_6 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  stage1_regs_r_0_0_7 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  stage1_regs_r_0_0_8 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  stage1_regs_r_0_1_0 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  stage1_regs_r_0_1_1 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  stage1_regs_r_0_1_2 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  stage1_regs_r_0_1_3 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  stage1_regs_r_0_1_4 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  stage1_regs_r_0_1_5 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  stage1_regs_r_0_1_6 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  stage1_regs_r_0_1_7 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  stage1_regs_r_0_1_8 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  stage1_regs_r_1_0_0 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  stage1_regs_r_1_0_1 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  stage1_regs_r_1_0_2 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  stage1_regs_r_1_0_3 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  stage1_regs_r_1_0_4 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  stage1_regs_r_1_0_5 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  stage1_regs_r_1_0_6 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  stage1_regs_r_1_0_7 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  stage1_regs_r_1_0_8 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  stage1_regs_r_1_1_0 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  stage1_regs_r_1_1_1 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  stage1_regs_r_1_1_2 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  stage1_regs_r_1_1_3 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  stage1_regs_r_1_1_4 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  stage1_regs_r_1_1_5 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  stage1_regs_r_1_1_6 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  stage1_regs_r_1_1_7 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_regs_r_1_1_8 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  stage2_regs_r_0_0_0 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  stage2_regs_r_0_0_1 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  stage2_regs_r_0_0_2 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  stage2_regs_r_0_0_3 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  stage2_regs_r_0_0_4 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  stage2_regs_r_0_0_5 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  stage2_regs_r_0_0_6 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  stage2_regs_r_0_0_7 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  stage2_regs_r_0_0_8 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  stage2_regs_r_0_0_9 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  stage2_regs_r_0_0_10 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  stage2_regs_r_0_0_11 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  stage2_regs_r_0_1_0 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  stage2_regs_r_0_1_1 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  stage2_regs_r_0_1_2 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  stage2_regs_r_0_1_3 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  stage2_regs_r_0_1_4 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  stage2_regs_r_0_1_5 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  stage2_regs_r_0_1_6 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  stage2_regs_r_0_1_7 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  stage2_regs_r_0_1_8 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  stage2_regs_r_0_1_9 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  stage2_regs_r_0_1_10 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  stage2_regs_r_0_1_11 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  stage2_regs_r_1_0_0 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  stage2_regs_r_1_0_1 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  stage2_regs_r_1_0_2 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  stage2_regs_r_1_0_3 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  stage2_regs_r_1_0_4 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  stage2_regs_r_1_0_5 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  stage2_regs_r_1_0_6 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  stage2_regs_r_1_0_7 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  stage2_regs_r_1_0_8 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  stage2_regs_r_1_0_9 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  stage2_regs_r_1_0_10 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  stage2_regs_r_1_0_11 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  stage2_regs_r_1_1_0 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  stage2_regs_r_1_1_1 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  stage2_regs_r_1_1_2 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  stage2_regs_r_1_1_3 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  stage2_regs_r_1_1_4 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  stage2_regs_r_1_1_5 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  stage2_regs_r_1_1_6 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  stage2_regs_r_1_1_7 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  stage2_regs_r_1_1_8 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  stage2_regs_r_1_1_9 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  stage2_regs_r_1_1_10 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  stage2_regs_r_1_1_11 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  stage3_regs_r_0_1_0 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  stage3_regs_r_0_1_1 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  stage3_regs_r_0_1_2 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  stage3_regs_r_0_1_3 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  stage3_regs_r_0_1_4 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  stage3_regs_r_0_1_5 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  stage3_regs_r_0_1_6 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  stage3_regs_r_0_1_7 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  stage3_regs_r_0_1_8 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  stage3_regs_r_1_1_0 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  stage3_regs_r_1_1_1 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  stage3_regs_r_1_1_2 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  stage3_regs_r_1_1_3 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  stage3_regs_r_1_1_4 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  stage3_regs_r_1_1_5 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  stage3_regs_r_1_1_6 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  stage3_regs_r_1_1_7 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  stage3_regs_r_1_1_8 = _RAND_197[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hqr7(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  output [31:0] io_out_s
);
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2533:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2533:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2533:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2533:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2533:28]
  wire  FP_reciprocal_newfpu_clock; // @[FloatingPointDesigns.scala 2534:28]
  wire  FP_reciprocal_newfpu_reset; // @[FloatingPointDesigns.scala 2534:28]
  wire [31:0] FP_reciprocal_newfpu_io_in_a; // @[FloatingPointDesigns.scala 2534:28]
  wire [31:0] FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2534:28]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2533:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_reciprocal_newfpu FP_reciprocal_newfpu ( // @[FloatingPointDesigns.scala 2534:28]
    .clock(FP_reciprocal_newfpu_clock),
    .reset(FP_reciprocal_newfpu_reset),
    .io_in_a(FP_reciprocal_newfpu_io_in_a),
    .io_out_s(FP_reciprocal_newfpu_io_out_s)
  );
  assign io_out_s = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2541:14]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = 32'hc0000000; // @[FloatingPointDesigns.scala 2538:21]
  assign FP_multiplier_10ccs_io_in_b = FP_reciprocal_newfpu_io_out_s; // @[FloatingPointDesigns.scala 2539:21]
  assign FP_reciprocal_newfpu_clock = clock;
  assign FP_reciprocal_newfpu_reset = reset;
  assign FP_reciprocal_newfpu_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2537:21]
endmodule
module FPReg(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] reg_0; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_1; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_2; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_3; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_4; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_5; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_6; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_7; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_8; // @[FloatingPointDesigns.scala 2270:22]
  reg [31:0] reg_9; // @[FloatingPointDesigns.scala 2270:22]
  assign io_out = reg_9; // @[FloatingPointDesigns.scala 2276:12]
  always @(posedge clock) begin
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_0 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_0 <= io_in; // @[FloatingPointDesigns.scala 2272:14]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_1 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_1 <= reg_0; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_2 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_2 <= reg_1; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_3 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_3 <= reg_2; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_4 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_4 <= reg_3; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_5 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_5 <= reg_4; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_6 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_6 <= reg_5; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_7 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_7 <= reg_6; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_8 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_8 <= reg_7; // @[FloatingPointDesigns.scala 2274:16]
    end
    if (reset) begin // @[FloatingPointDesigns.scala 2270:22]
      reg_9 <= 32'h0; // @[FloatingPointDesigns.scala 2270:22]
    end else begin
      reg_9 <= reg_8; // @[FloatingPointDesigns.scala 2274:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_9 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axpy_dp(
  input         clock,
  input         reset,
  input  [31:0] io_in_a,
  input  [31:0] io_in_b_0,
  input  [31:0] io_in_b_1,
  input  [31:0] io_in_b_2,
  input  [31:0] io_in_b_3,
  input  [31:0] io_in_b_4,
  input  [31:0] io_in_b_5,
  input  [31:0] io_in_b_6,
  input  [31:0] io_in_b_7,
  input  [31:0] io_in_b_8,
  input  [31:0] io_in_b_9,
  input  [31:0] io_in_b_10,
  input  [31:0] io_in_b_11,
  input  [31:0] io_in_b_12,
  input  [31:0] io_in_b_13,
  input  [31:0] io_in_b_14,
  input  [31:0] io_in_b_15,
  input  [31:0] io_in_b_16,
  input  [31:0] io_in_b_17,
  input  [31:0] io_in_b_18,
  input  [31:0] io_in_b_19,
  input  [31:0] io_in_b_20,
  input  [31:0] io_in_b_21,
  input  [31:0] io_in_b_22,
  input  [31:0] io_in_b_23,
  input  [31:0] io_in_b_24,
  input  [31:0] io_in_b_25,
  input  [31:0] io_in_b_26,
  input  [31:0] io_in_b_27,
  input  [31:0] io_in_b_28,
  input  [31:0] io_in_b_29,
  input  [31:0] io_in_b_30,
  input  [31:0] io_in_b_31,
  input  [31:0] io_in_b_32,
  input  [31:0] io_in_b_33,
  input  [31:0] io_in_b_34,
  input  [31:0] io_in_b_35,
  input  [31:0] io_in_b_36,
  input  [31:0] io_in_b_37,
  input  [31:0] io_in_b_38,
  input  [31:0] io_in_b_39,
  input  [31:0] io_in_b_40,
  input  [31:0] io_in_b_41,
  input  [31:0] io_in_b_42,
  input  [31:0] io_in_b_43,
  input  [31:0] io_in_b_44,
  input  [31:0] io_in_b_45,
  input  [31:0] io_in_b_46,
  input  [31:0] io_in_b_47,
  input  [31:0] io_in_b_48,
  input  [31:0] io_in_b_49,
  input  [31:0] io_in_b_50,
  input  [31:0] io_in_b_51,
  input  [31:0] io_in_b_52,
  input  [31:0] io_in_b_53,
  input  [31:0] io_in_b_54,
  input  [31:0] io_in_b_55,
  input  [31:0] io_in_b_56,
  input  [31:0] io_in_b_57,
  input  [31:0] io_in_b_58,
  input  [31:0] io_in_b_59,
  input  [31:0] io_in_b_60,
  input  [31:0] io_in_b_61,
  input  [31:0] io_in_b_62,
  input  [31:0] io_in_b_63,
  input  [31:0] io_in_c_0,
  input  [31:0] io_in_c_1,
  input  [31:0] io_in_c_2,
  input  [31:0] io_in_c_3,
  input  [31:0] io_in_c_4,
  input  [31:0] io_in_c_5,
  input  [31:0] io_in_c_6,
  input  [31:0] io_in_c_7,
  input  [31:0] io_in_c_8,
  input  [31:0] io_in_c_9,
  input  [31:0] io_in_c_10,
  input  [31:0] io_in_c_11,
  input  [31:0] io_in_c_12,
  input  [31:0] io_in_c_13,
  input  [31:0] io_in_c_14,
  input  [31:0] io_in_c_15,
  input  [31:0] io_in_c_16,
  input  [31:0] io_in_c_17,
  input  [31:0] io_in_c_18,
  input  [31:0] io_in_c_19,
  input  [31:0] io_in_c_20,
  input  [31:0] io_in_c_21,
  input  [31:0] io_in_c_22,
  input  [31:0] io_in_c_23,
  input  [31:0] io_in_c_24,
  input  [31:0] io_in_c_25,
  input  [31:0] io_in_c_26,
  input  [31:0] io_in_c_27,
  input  [31:0] io_in_c_28,
  input  [31:0] io_in_c_29,
  input  [31:0] io_in_c_30,
  input  [31:0] io_in_c_31,
  input  [31:0] io_in_c_32,
  input  [31:0] io_in_c_33,
  input  [31:0] io_in_c_34,
  input  [31:0] io_in_c_35,
  input  [31:0] io_in_c_36,
  input  [31:0] io_in_c_37,
  input  [31:0] io_in_c_38,
  input  [31:0] io_in_c_39,
  input  [31:0] io_in_c_40,
  input  [31:0] io_in_c_41,
  input  [31:0] io_in_c_42,
  input  [31:0] io_in_c_43,
  input  [31:0] io_in_c_44,
  input  [31:0] io_in_c_45,
  input  [31:0] io_in_c_46,
  input  [31:0] io_in_c_47,
  input  [31:0] io_in_c_48,
  input  [31:0] io_in_c_49,
  input  [31:0] io_in_c_50,
  input  [31:0] io_in_c_51,
  input  [31:0] io_in_c_52,
  input  [31:0] io_in_c_53,
  input  [31:0] io_in_c_54,
  input  [31:0] io_in_c_55,
  input  [31:0] io_in_c_56,
  input  [31:0] io_in_c_57,
  input  [31:0] io_in_c_58,
  input  [31:0] io_in_c_59,
  input  [31:0] io_in_c_60,
  input  [31:0] io_in_c_61,
  input  [31:0] io_in_c_62,
  input  [31:0] io_in_c_63,
  output [31:0] io_out_s_0,
  output [31:0] io_out_s_1,
  output [31:0] io_out_s_2,
  output [31:0] io_out_s_3,
  output [31:0] io_out_s_4,
  output [31:0] io_out_s_5,
  output [31:0] io_out_s_6,
  output [31:0] io_out_s_7,
  output [31:0] io_out_s_8,
  output [31:0] io_out_s_9,
  output [31:0] io_out_s_10,
  output [31:0] io_out_s_11,
  output [31:0] io_out_s_12,
  output [31:0] io_out_s_13,
  output [31:0] io_out_s_14,
  output [31:0] io_out_s_15,
  output [31:0] io_out_s_16,
  output [31:0] io_out_s_17,
  output [31:0] io_out_s_18,
  output [31:0] io_out_s_19,
  output [31:0] io_out_s_20,
  output [31:0] io_out_s_21,
  output [31:0] io_out_s_22,
  output [31:0] io_out_s_23,
  output [31:0] io_out_s_24,
  output [31:0] io_out_s_25,
  output [31:0] io_out_s_26,
  output [31:0] io_out_s_27,
  output [31:0] io_out_s_28,
  output [31:0] io_out_s_29,
  output [31:0] io_out_s_30,
  output [31:0] io_out_s_31,
  output [31:0] io_out_s_32,
  output [31:0] io_out_s_33,
  output [31:0] io_out_s_34,
  output [31:0] io_out_s_35,
  output [31:0] io_out_s_36,
  output [31:0] io_out_s_37,
  output [31:0] io_out_s_38,
  output [31:0] io_out_s_39,
  output [31:0] io_out_s_40,
  output [31:0] io_out_s_41,
  output [31:0] io_out_s_42,
  output [31:0] io_out_s_43,
  output [31:0] io_out_s_44,
  output [31:0] io_out_s_45,
  output [31:0] io_out_s_46,
  output [31:0] io_out_s_47,
  output [31:0] io_out_s_48,
  output [31:0] io_out_s_49,
  output [31:0] io_out_s_50,
  output [31:0] io_out_s_51,
  output [31:0] io_out_s_52,
  output [31:0] io_out_s_53,
  output [31:0] io_out_s_54,
  output [31:0] io_out_s_55,
  output [31:0] io_out_s_56,
  output [31:0] io_out_s_57,
  output [31:0] io_out_s_58,
  output [31:0] io_out_s_59,
  output [31:0] io_out_s_60,
  output [31:0] io_out_s_61,
  output [31:0] io_out_s_62,
  output [31:0] io_out_s_63
);
  wire  FP_multiplier_10ccs_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_1_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_1_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_2_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_2_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_3_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_3_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_4_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_4_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_5_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_5_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_6_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_6_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_7_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_7_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_8_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_8_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_9_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_9_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_10_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_10_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_11_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_11_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_12_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_12_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_13_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_13_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_14_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_14_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_15_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_15_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_16_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_16_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_17_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_17_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_18_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_18_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_19_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_19_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_20_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_20_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_21_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_21_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_22_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_22_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_23_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_23_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_24_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_24_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_25_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_25_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_26_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_26_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_27_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_27_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_28_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_28_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_29_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_29_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_30_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_30_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_31_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_31_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_32_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_32_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_33_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_33_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_34_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_34_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_35_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_35_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_36_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_36_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_37_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_37_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_38_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_38_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_39_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_39_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_40_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_40_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_41_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_41_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_42_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_42_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_43_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_43_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_44_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_44_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_45_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_45_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_46_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_46_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_47_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_47_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_48_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_48_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_49_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_49_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_50_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_50_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_51_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_51_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_52_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_52_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_53_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_53_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_54_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_54_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_55_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_55_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_56_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_56_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_57_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_57_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_58_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_58_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_59_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_59_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_60_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_60_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_61_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_61_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_62_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_62_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_63_clock; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_multiplier_10ccs_63_reset; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2485:28]
  wire [31:0] FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2485:28]
  wire  FP_adder_13ccs_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_1_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_1_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_1_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_1_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_2_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_2_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_2_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_2_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_3_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_3_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_3_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_3_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_4_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_4_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_4_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_4_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_5_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_5_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_5_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_5_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_6_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_6_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_6_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_6_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_7_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_7_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_7_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_7_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_8_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_8_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_8_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_8_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_9_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_9_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_9_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_9_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_10_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_10_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_10_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_10_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_11_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_11_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_11_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_11_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_12_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_12_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_12_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_12_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_13_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_13_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_13_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_13_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_14_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_14_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_14_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_14_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_15_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_15_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_15_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_15_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_16_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_16_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_16_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_16_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_17_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_17_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_17_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_17_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_18_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_18_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_18_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_18_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_19_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_19_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_19_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_19_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_20_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_20_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_20_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_20_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_21_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_21_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_21_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_21_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_22_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_22_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_22_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_22_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_23_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_23_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_23_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_23_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_24_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_24_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_24_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_24_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_25_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_25_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_25_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_25_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_26_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_26_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_26_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_26_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_27_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_27_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_27_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_27_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_28_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_28_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_28_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_28_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_29_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_29_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_29_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_29_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_30_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_30_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_30_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_30_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_31_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_31_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_31_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_31_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_32_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_32_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_32_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_32_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_33_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_33_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_33_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_33_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_34_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_34_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_34_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_34_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_35_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_35_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_35_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_35_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_36_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_36_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_36_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_36_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_37_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_37_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_37_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_37_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_38_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_38_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_38_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_38_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_39_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_39_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_39_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_39_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_40_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_40_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_40_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_40_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_41_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_41_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_41_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_41_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_42_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_42_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_42_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_42_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_43_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_43_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_43_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_43_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_44_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_44_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_44_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_44_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_45_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_45_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_45_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_45_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_46_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_46_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_46_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_46_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_47_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_47_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_47_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_47_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_48_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_48_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_48_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_48_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_49_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_49_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_49_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_49_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_50_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_50_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_50_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_50_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_51_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_51_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_51_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_51_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_52_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_52_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_52_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_52_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_53_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_53_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_53_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_53_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_54_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_54_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_54_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_54_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_55_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_55_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_55_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_55_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_56_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_56_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_56_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_56_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_57_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_57_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_57_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_57_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_58_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_58_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_58_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_58_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_59_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_59_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_59_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_59_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_60_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_60_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_60_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_60_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_61_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_61_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_61_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_61_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_62_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_62_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_62_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_62_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_63_clock; // @[FloatingPointDesigns.scala 2490:25]
  wire  FP_adder_13ccs_63_reset; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_63_io_in_a; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_63_io_in_b; // @[FloatingPointDesigns.scala 2490:25]
  wire [31:0] FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2490:25]
  wire  FPReg_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_1_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_1_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_1_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_1_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_2_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_2_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_2_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_2_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_3_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_3_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_3_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_3_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_4_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_4_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_4_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_4_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_5_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_5_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_5_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_5_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_6_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_6_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_6_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_6_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_7_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_7_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_7_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_7_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_8_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_8_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_8_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_8_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_9_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_9_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_9_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_9_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_10_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_10_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_10_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_10_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_11_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_11_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_11_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_11_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_12_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_12_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_12_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_12_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_13_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_13_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_13_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_13_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_14_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_14_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_14_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_14_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_15_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_15_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_15_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_15_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_16_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_16_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_16_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_16_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_17_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_17_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_17_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_17_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_18_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_18_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_18_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_18_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_19_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_19_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_19_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_19_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_20_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_20_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_20_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_20_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_21_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_21_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_21_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_21_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_22_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_22_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_22_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_22_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_23_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_23_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_23_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_23_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_24_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_24_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_24_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_24_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_25_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_25_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_25_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_25_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_26_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_26_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_26_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_26_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_27_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_27_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_27_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_27_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_28_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_28_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_28_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_28_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_29_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_29_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_29_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_29_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_30_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_30_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_30_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_30_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_31_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_31_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_31_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_31_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_32_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_32_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_32_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_32_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_33_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_33_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_33_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_33_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_34_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_34_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_34_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_34_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_35_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_35_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_35_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_35_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_36_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_36_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_36_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_36_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_37_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_37_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_37_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_37_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_38_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_38_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_38_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_38_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_39_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_39_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_39_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_39_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_40_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_40_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_40_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_40_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_41_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_41_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_41_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_41_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_42_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_42_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_42_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_42_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_43_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_43_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_43_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_43_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_44_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_44_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_44_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_44_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_45_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_45_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_45_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_45_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_46_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_46_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_46_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_46_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_47_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_47_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_47_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_47_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_48_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_48_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_48_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_48_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_49_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_49_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_49_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_49_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_50_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_50_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_50_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_50_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_51_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_51_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_51_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_51_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_52_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_52_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_52_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_52_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_53_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_53_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_53_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_53_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_54_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_54_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_54_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_54_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_55_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_55_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_55_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_55_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_56_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_56_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_56_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_56_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_57_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_57_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_57_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_57_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_58_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_58_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_58_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_58_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_59_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_59_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_59_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_59_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_60_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_60_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_60_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_60_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_61_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_61_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_61_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_61_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_62_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_62_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_62_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_62_io_out; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_63_clock; // @[FloatingPointDesigns.scala 2494:48]
  wire  FPReg_63_reset; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_63_io_in; // @[FloatingPointDesigns.scala 2494:48]
  wire [31:0] FPReg_63_io_out; // @[FloatingPointDesigns.scala 2494:48]
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_1 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_1_clock),
    .reset(FP_multiplier_10ccs_1_reset),
    .io_in_a(FP_multiplier_10ccs_1_io_in_a),
    .io_in_b(FP_multiplier_10ccs_1_io_in_b),
    .io_out_s(FP_multiplier_10ccs_1_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_2 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_2_clock),
    .reset(FP_multiplier_10ccs_2_reset),
    .io_in_a(FP_multiplier_10ccs_2_io_in_a),
    .io_in_b(FP_multiplier_10ccs_2_io_in_b),
    .io_out_s(FP_multiplier_10ccs_2_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_3 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_3_clock),
    .reset(FP_multiplier_10ccs_3_reset),
    .io_in_a(FP_multiplier_10ccs_3_io_in_a),
    .io_in_b(FP_multiplier_10ccs_3_io_in_b),
    .io_out_s(FP_multiplier_10ccs_3_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_4 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_4_clock),
    .reset(FP_multiplier_10ccs_4_reset),
    .io_in_a(FP_multiplier_10ccs_4_io_in_a),
    .io_in_b(FP_multiplier_10ccs_4_io_in_b),
    .io_out_s(FP_multiplier_10ccs_4_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_5 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_5_clock),
    .reset(FP_multiplier_10ccs_5_reset),
    .io_in_a(FP_multiplier_10ccs_5_io_in_a),
    .io_in_b(FP_multiplier_10ccs_5_io_in_b),
    .io_out_s(FP_multiplier_10ccs_5_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_6 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_6_clock),
    .reset(FP_multiplier_10ccs_6_reset),
    .io_in_a(FP_multiplier_10ccs_6_io_in_a),
    .io_in_b(FP_multiplier_10ccs_6_io_in_b),
    .io_out_s(FP_multiplier_10ccs_6_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_7 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_7_clock),
    .reset(FP_multiplier_10ccs_7_reset),
    .io_in_a(FP_multiplier_10ccs_7_io_in_a),
    .io_in_b(FP_multiplier_10ccs_7_io_in_b),
    .io_out_s(FP_multiplier_10ccs_7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_8 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_8_clock),
    .reset(FP_multiplier_10ccs_8_reset),
    .io_in_a(FP_multiplier_10ccs_8_io_in_a),
    .io_in_b(FP_multiplier_10ccs_8_io_in_b),
    .io_out_s(FP_multiplier_10ccs_8_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_9 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_9_clock),
    .reset(FP_multiplier_10ccs_9_reset),
    .io_in_a(FP_multiplier_10ccs_9_io_in_a),
    .io_in_b(FP_multiplier_10ccs_9_io_in_b),
    .io_out_s(FP_multiplier_10ccs_9_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_10 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_10_clock),
    .reset(FP_multiplier_10ccs_10_reset),
    .io_in_a(FP_multiplier_10ccs_10_io_in_a),
    .io_in_b(FP_multiplier_10ccs_10_io_in_b),
    .io_out_s(FP_multiplier_10ccs_10_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_11 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_11_clock),
    .reset(FP_multiplier_10ccs_11_reset),
    .io_in_a(FP_multiplier_10ccs_11_io_in_a),
    .io_in_b(FP_multiplier_10ccs_11_io_in_b),
    .io_out_s(FP_multiplier_10ccs_11_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_12 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_12_clock),
    .reset(FP_multiplier_10ccs_12_reset),
    .io_in_a(FP_multiplier_10ccs_12_io_in_a),
    .io_in_b(FP_multiplier_10ccs_12_io_in_b),
    .io_out_s(FP_multiplier_10ccs_12_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_13 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_13_clock),
    .reset(FP_multiplier_10ccs_13_reset),
    .io_in_a(FP_multiplier_10ccs_13_io_in_a),
    .io_in_b(FP_multiplier_10ccs_13_io_in_b),
    .io_out_s(FP_multiplier_10ccs_13_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_14 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_14_clock),
    .reset(FP_multiplier_10ccs_14_reset),
    .io_in_a(FP_multiplier_10ccs_14_io_in_a),
    .io_in_b(FP_multiplier_10ccs_14_io_in_b),
    .io_out_s(FP_multiplier_10ccs_14_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_15 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_15_clock),
    .reset(FP_multiplier_10ccs_15_reset),
    .io_in_a(FP_multiplier_10ccs_15_io_in_a),
    .io_in_b(FP_multiplier_10ccs_15_io_in_b),
    .io_out_s(FP_multiplier_10ccs_15_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_16 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_16_clock),
    .reset(FP_multiplier_10ccs_16_reset),
    .io_in_a(FP_multiplier_10ccs_16_io_in_a),
    .io_in_b(FP_multiplier_10ccs_16_io_in_b),
    .io_out_s(FP_multiplier_10ccs_16_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_17 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_17_clock),
    .reset(FP_multiplier_10ccs_17_reset),
    .io_in_a(FP_multiplier_10ccs_17_io_in_a),
    .io_in_b(FP_multiplier_10ccs_17_io_in_b),
    .io_out_s(FP_multiplier_10ccs_17_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_18 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_18_clock),
    .reset(FP_multiplier_10ccs_18_reset),
    .io_in_a(FP_multiplier_10ccs_18_io_in_a),
    .io_in_b(FP_multiplier_10ccs_18_io_in_b),
    .io_out_s(FP_multiplier_10ccs_18_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_19 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_19_clock),
    .reset(FP_multiplier_10ccs_19_reset),
    .io_in_a(FP_multiplier_10ccs_19_io_in_a),
    .io_in_b(FP_multiplier_10ccs_19_io_in_b),
    .io_out_s(FP_multiplier_10ccs_19_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_20 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_20_clock),
    .reset(FP_multiplier_10ccs_20_reset),
    .io_in_a(FP_multiplier_10ccs_20_io_in_a),
    .io_in_b(FP_multiplier_10ccs_20_io_in_b),
    .io_out_s(FP_multiplier_10ccs_20_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_21 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_21_clock),
    .reset(FP_multiplier_10ccs_21_reset),
    .io_in_a(FP_multiplier_10ccs_21_io_in_a),
    .io_in_b(FP_multiplier_10ccs_21_io_in_b),
    .io_out_s(FP_multiplier_10ccs_21_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_22 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_22_clock),
    .reset(FP_multiplier_10ccs_22_reset),
    .io_in_a(FP_multiplier_10ccs_22_io_in_a),
    .io_in_b(FP_multiplier_10ccs_22_io_in_b),
    .io_out_s(FP_multiplier_10ccs_22_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_23 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_23_clock),
    .reset(FP_multiplier_10ccs_23_reset),
    .io_in_a(FP_multiplier_10ccs_23_io_in_a),
    .io_in_b(FP_multiplier_10ccs_23_io_in_b),
    .io_out_s(FP_multiplier_10ccs_23_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_24 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_24_clock),
    .reset(FP_multiplier_10ccs_24_reset),
    .io_in_a(FP_multiplier_10ccs_24_io_in_a),
    .io_in_b(FP_multiplier_10ccs_24_io_in_b),
    .io_out_s(FP_multiplier_10ccs_24_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_25 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_25_clock),
    .reset(FP_multiplier_10ccs_25_reset),
    .io_in_a(FP_multiplier_10ccs_25_io_in_a),
    .io_in_b(FP_multiplier_10ccs_25_io_in_b),
    .io_out_s(FP_multiplier_10ccs_25_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_26 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_26_clock),
    .reset(FP_multiplier_10ccs_26_reset),
    .io_in_a(FP_multiplier_10ccs_26_io_in_a),
    .io_in_b(FP_multiplier_10ccs_26_io_in_b),
    .io_out_s(FP_multiplier_10ccs_26_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_27 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_27_clock),
    .reset(FP_multiplier_10ccs_27_reset),
    .io_in_a(FP_multiplier_10ccs_27_io_in_a),
    .io_in_b(FP_multiplier_10ccs_27_io_in_b),
    .io_out_s(FP_multiplier_10ccs_27_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_28 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_28_clock),
    .reset(FP_multiplier_10ccs_28_reset),
    .io_in_a(FP_multiplier_10ccs_28_io_in_a),
    .io_in_b(FP_multiplier_10ccs_28_io_in_b),
    .io_out_s(FP_multiplier_10ccs_28_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_29 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_29_clock),
    .reset(FP_multiplier_10ccs_29_reset),
    .io_in_a(FP_multiplier_10ccs_29_io_in_a),
    .io_in_b(FP_multiplier_10ccs_29_io_in_b),
    .io_out_s(FP_multiplier_10ccs_29_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_30 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_30_clock),
    .reset(FP_multiplier_10ccs_30_reset),
    .io_in_a(FP_multiplier_10ccs_30_io_in_a),
    .io_in_b(FP_multiplier_10ccs_30_io_in_b),
    .io_out_s(FP_multiplier_10ccs_30_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_31 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_31_clock),
    .reset(FP_multiplier_10ccs_31_reset),
    .io_in_a(FP_multiplier_10ccs_31_io_in_a),
    .io_in_b(FP_multiplier_10ccs_31_io_in_b),
    .io_out_s(FP_multiplier_10ccs_31_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_32 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_32_clock),
    .reset(FP_multiplier_10ccs_32_reset),
    .io_in_a(FP_multiplier_10ccs_32_io_in_a),
    .io_in_b(FP_multiplier_10ccs_32_io_in_b),
    .io_out_s(FP_multiplier_10ccs_32_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_33 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_33_clock),
    .reset(FP_multiplier_10ccs_33_reset),
    .io_in_a(FP_multiplier_10ccs_33_io_in_a),
    .io_in_b(FP_multiplier_10ccs_33_io_in_b),
    .io_out_s(FP_multiplier_10ccs_33_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_34 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_34_clock),
    .reset(FP_multiplier_10ccs_34_reset),
    .io_in_a(FP_multiplier_10ccs_34_io_in_a),
    .io_in_b(FP_multiplier_10ccs_34_io_in_b),
    .io_out_s(FP_multiplier_10ccs_34_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_35 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_35_clock),
    .reset(FP_multiplier_10ccs_35_reset),
    .io_in_a(FP_multiplier_10ccs_35_io_in_a),
    .io_in_b(FP_multiplier_10ccs_35_io_in_b),
    .io_out_s(FP_multiplier_10ccs_35_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_36 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_36_clock),
    .reset(FP_multiplier_10ccs_36_reset),
    .io_in_a(FP_multiplier_10ccs_36_io_in_a),
    .io_in_b(FP_multiplier_10ccs_36_io_in_b),
    .io_out_s(FP_multiplier_10ccs_36_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_37 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_37_clock),
    .reset(FP_multiplier_10ccs_37_reset),
    .io_in_a(FP_multiplier_10ccs_37_io_in_a),
    .io_in_b(FP_multiplier_10ccs_37_io_in_b),
    .io_out_s(FP_multiplier_10ccs_37_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_38 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_38_clock),
    .reset(FP_multiplier_10ccs_38_reset),
    .io_in_a(FP_multiplier_10ccs_38_io_in_a),
    .io_in_b(FP_multiplier_10ccs_38_io_in_b),
    .io_out_s(FP_multiplier_10ccs_38_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_39 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_39_clock),
    .reset(FP_multiplier_10ccs_39_reset),
    .io_in_a(FP_multiplier_10ccs_39_io_in_a),
    .io_in_b(FP_multiplier_10ccs_39_io_in_b),
    .io_out_s(FP_multiplier_10ccs_39_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_40 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_40_clock),
    .reset(FP_multiplier_10ccs_40_reset),
    .io_in_a(FP_multiplier_10ccs_40_io_in_a),
    .io_in_b(FP_multiplier_10ccs_40_io_in_b),
    .io_out_s(FP_multiplier_10ccs_40_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_41 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_41_clock),
    .reset(FP_multiplier_10ccs_41_reset),
    .io_in_a(FP_multiplier_10ccs_41_io_in_a),
    .io_in_b(FP_multiplier_10ccs_41_io_in_b),
    .io_out_s(FP_multiplier_10ccs_41_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_42 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_42_clock),
    .reset(FP_multiplier_10ccs_42_reset),
    .io_in_a(FP_multiplier_10ccs_42_io_in_a),
    .io_in_b(FP_multiplier_10ccs_42_io_in_b),
    .io_out_s(FP_multiplier_10ccs_42_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_43 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_43_clock),
    .reset(FP_multiplier_10ccs_43_reset),
    .io_in_a(FP_multiplier_10ccs_43_io_in_a),
    .io_in_b(FP_multiplier_10ccs_43_io_in_b),
    .io_out_s(FP_multiplier_10ccs_43_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_44 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_44_clock),
    .reset(FP_multiplier_10ccs_44_reset),
    .io_in_a(FP_multiplier_10ccs_44_io_in_a),
    .io_in_b(FP_multiplier_10ccs_44_io_in_b),
    .io_out_s(FP_multiplier_10ccs_44_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_45 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_45_clock),
    .reset(FP_multiplier_10ccs_45_reset),
    .io_in_a(FP_multiplier_10ccs_45_io_in_a),
    .io_in_b(FP_multiplier_10ccs_45_io_in_b),
    .io_out_s(FP_multiplier_10ccs_45_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_46 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_46_clock),
    .reset(FP_multiplier_10ccs_46_reset),
    .io_in_a(FP_multiplier_10ccs_46_io_in_a),
    .io_in_b(FP_multiplier_10ccs_46_io_in_b),
    .io_out_s(FP_multiplier_10ccs_46_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_47 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_47_clock),
    .reset(FP_multiplier_10ccs_47_reset),
    .io_in_a(FP_multiplier_10ccs_47_io_in_a),
    .io_in_b(FP_multiplier_10ccs_47_io_in_b),
    .io_out_s(FP_multiplier_10ccs_47_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_48 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_48_clock),
    .reset(FP_multiplier_10ccs_48_reset),
    .io_in_a(FP_multiplier_10ccs_48_io_in_a),
    .io_in_b(FP_multiplier_10ccs_48_io_in_b),
    .io_out_s(FP_multiplier_10ccs_48_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_49 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_49_clock),
    .reset(FP_multiplier_10ccs_49_reset),
    .io_in_a(FP_multiplier_10ccs_49_io_in_a),
    .io_in_b(FP_multiplier_10ccs_49_io_in_b),
    .io_out_s(FP_multiplier_10ccs_49_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_50 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_50_clock),
    .reset(FP_multiplier_10ccs_50_reset),
    .io_in_a(FP_multiplier_10ccs_50_io_in_a),
    .io_in_b(FP_multiplier_10ccs_50_io_in_b),
    .io_out_s(FP_multiplier_10ccs_50_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_51 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_51_clock),
    .reset(FP_multiplier_10ccs_51_reset),
    .io_in_a(FP_multiplier_10ccs_51_io_in_a),
    .io_in_b(FP_multiplier_10ccs_51_io_in_b),
    .io_out_s(FP_multiplier_10ccs_51_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_52 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_52_clock),
    .reset(FP_multiplier_10ccs_52_reset),
    .io_in_a(FP_multiplier_10ccs_52_io_in_a),
    .io_in_b(FP_multiplier_10ccs_52_io_in_b),
    .io_out_s(FP_multiplier_10ccs_52_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_53 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_53_clock),
    .reset(FP_multiplier_10ccs_53_reset),
    .io_in_a(FP_multiplier_10ccs_53_io_in_a),
    .io_in_b(FP_multiplier_10ccs_53_io_in_b),
    .io_out_s(FP_multiplier_10ccs_53_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_54 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_54_clock),
    .reset(FP_multiplier_10ccs_54_reset),
    .io_in_a(FP_multiplier_10ccs_54_io_in_a),
    .io_in_b(FP_multiplier_10ccs_54_io_in_b),
    .io_out_s(FP_multiplier_10ccs_54_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_55 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_55_clock),
    .reset(FP_multiplier_10ccs_55_reset),
    .io_in_a(FP_multiplier_10ccs_55_io_in_a),
    .io_in_b(FP_multiplier_10ccs_55_io_in_b),
    .io_out_s(FP_multiplier_10ccs_55_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_56 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_56_clock),
    .reset(FP_multiplier_10ccs_56_reset),
    .io_in_a(FP_multiplier_10ccs_56_io_in_a),
    .io_in_b(FP_multiplier_10ccs_56_io_in_b),
    .io_out_s(FP_multiplier_10ccs_56_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_57 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_57_clock),
    .reset(FP_multiplier_10ccs_57_reset),
    .io_in_a(FP_multiplier_10ccs_57_io_in_a),
    .io_in_b(FP_multiplier_10ccs_57_io_in_b),
    .io_out_s(FP_multiplier_10ccs_57_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_58 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_58_clock),
    .reset(FP_multiplier_10ccs_58_reset),
    .io_in_a(FP_multiplier_10ccs_58_io_in_a),
    .io_in_b(FP_multiplier_10ccs_58_io_in_b),
    .io_out_s(FP_multiplier_10ccs_58_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_59 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_59_clock),
    .reset(FP_multiplier_10ccs_59_reset),
    .io_in_a(FP_multiplier_10ccs_59_io_in_a),
    .io_in_b(FP_multiplier_10ccs_59_io_in_b),
    .io_out_s(FP_multiplier_10ccs_59_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_60 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_60_clock),
    .reset(FP_multiplier_10ccs_60_reset),
    .io_in_a(FP_multiplier_10ccs_60_io_in_a),
    .io_in_b(FP_multiplier_10ccs_60_io_in_b),
    .io_out_s(FP_multiplier_10ccs_60_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_61 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_61_clock),
    .reset(FP_multiplier_10ccs_61_reset),
    .io_in_a(FP_multiplier_10ccs_61_io_in_a),
    .io_in_b(FP_multiplier_10ccs_61_io_in_b),
    .io_out_s(FP_multiplier_10ccs_61_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_62 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_62_clock),
    .reset(FP_multiplier_10ccs_62_reset),
    .io_in_a(FP_multiplier_10ccs_62_io_in_a),
    .io_in_b(FP_multiplier_10ccs_62_io_in_b),
    .io_out_s(FP_multiplier_10ccs_62_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs_63 ( // @[FloatingPointDesigns.scala 2485:28]
    .clock(FP_multiplier_10ccs_63_clock),
    .reset(FP_multiplier_10ccs_63_reset),
    .io_in_a(FP_multiplier_10ccs_63_io_in_a),
    .io_in_b(FP_multiplier_10ccs_63_io_in_b),
    .io_out_s(FP_multiplier_10ccs_63_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_clock),
    .reset(FP_adder_13ccs_reset),
    .io_in_a(FP_adder_13ccs_io_in_a),
    .io_in_b(FP_adder_13ccs_io_in_b),
    .io_out_s(FP_adder_13ccs_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_1 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_1_clock),
    .reset(FP_adder_13ccs_1_reset),
    .io_in_a(FP_adder_13ccs_1_io_in_a),
    .io_in_b(FP_adder_13ccs_1_io_in_b),
    .io_out_s(FP_adder_13ccs_1_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_2 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_2_clock),
    .reset(FP_adder_13ccs_2_reset),
    .io_in_a(FP_adder_13ccs_2_io_in_a),
    .io_in_b(FP_adder_13ccs_2_io_in_b),
    .io_out_s(FP_adder_13ccs_2_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_3 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_3_clock),
    .reset(FP_adder_13ccs_3_reset),
    .io_in_a(FP_adder_13ccs_3_io_in_a),
    .io_in_b(FP_adder_13ccs_3_io_in_b),
    .io_out_s(FP_adder_13ccs_3_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_4 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_4_clock),
    .reset(FP_adder_13ccs_4_reset),
    .io_in_a(FP_adder_13ccs_4_io_in_a),
    .io_in_b(FP_adder_13ccs_4_io_in_b),
    .io_out_s(FP_adder_13ccs_4_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_5 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_5_clock),
    .reset(FP_adder_13ccs_5_reset),
    .io_in_a(FP_adder_13ccs_5_io_in_a),
    .io_in_b(FP_adder_13ccs_5_io_in_b),
    .io_out_s(FP_adder_13ccs_5_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_6 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_6_clock),
    .reset(FP_adder_13ccs_6_reset),
    .io_in_a(FP_adder_13ccs_6_io_in_a),
    .io_in_b(FP_adder_13ccs_6_io_in_b),
    .io_out_s(FP_adder_13ccs_6_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_7 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_7_clock),
    .reset(FP_adder_13ccs_7_reset),
    .io_in_a(FP_adder_13ccs_7_io_in_a),
    .io_in_b(FP_adder_13ccs_7_io_in_b),
    .io_out_s(FP_adder_13ccs_7_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_8 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_8_clock),
    .reset(FP_adder_13ccs_8_reset),
    .io_in_a(FP_adder_13ccs_8_io_in_a),
    .io_in_b(FP_adder_13ccs_8_io_in_b),
    .io_out_s(FP_adder_13ccs_8_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_9 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_9_clock),
    .reset(FP_adder_13ccs_9_reset),
    .io_in_a(FP_adder_13ccs_9_io_in_a),
    .io_in_b(FP_adder_13ccs_9_io_in_b),
    .io_out_s(FP_adder_13ccs_9_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_10 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_10_clock),
    .reset(FP_adder_13ccs_10_reset),
    .io_in_a(FP_adder_13ccs_10_io_in_a),
    .io_in_b(FP_adder_13ccs_10_io_in_b),
    .io_out_s(FP_adder_13ccs_10_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_11 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_11_clock),
    .reset(FP_adder_13ccs_11_reset),
    .io_in_a(FP_adder_13ccs_11_io_in_a),
    .io_in_b(FP_adder_13ccs_11_io_in_b),
    .io_out_s(FP_adder_13ccs_11_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_12 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_12_clock),
    .reset(FP_adder_13ccs_12_reset),
    .io_in_a(FP_adder_13ccs_12_io_in_a),
    .io_in_b(FP_adder_13ccs_12_io_in_b),
    .io_out_s(FP_adder_13ccs_12_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_13 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_13_clock),
    .reset(FP_adder_13ccs_13_reset),
    .io_in_a(FP_adder_13ccs_13_io_in_a),
    .io_in_b(FP_adder_13ccs_13_io_in_b),
    .io_out_s(FP_adder_13ccs_13_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_14 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_14_clock),
    .reset(FP_adder_13ccs_14_reset),
    .io_in_a(FP_adder_13ccs_14_io_in_a),
    .io_in_b(FP_adder_13ccs_14_io_in_b),
    .io_out_s(FP_adder_13ccs_14_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_15 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_15_clock),
    .reset(FP_adder_13ccs_15_reset),
    .io_in_a(FP_adder_13ccs_15_io_in_a),
    .io_in_b(FP_adder_13ccs_15_io_in_b),
    .io_out_s(FP_adder_13ccs_15_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_16 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_16_clock),
    .reset(FP_adder_13ccs_16_reset),
    .io_in_a(FP_adder_13ccs_16_io_in_a),
    .io_in_b(FP_adder_13ccs_16_io_in_b),
    .io_out_s(FP_adder_13ccs_16_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_17 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_17_clock),
    .reset(FP_adder_13ccs_17_reset),
    .io_in_a(FP_adder_13ccs_17_io_in_a),
    .io_in_b(FP_adder_13ccs_17_io_in_b),
    .io_out_s(FP_adder_13ccs_17_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_18 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_18_clock),
    .reset(FP_adder_13ccs_18_reset),
    .io_in_a(FP_adder_13ccs_18_io_in_a),
    .io_in_b(FP_adder_13ccs_18_io_in_b),
    .io_out_s(FP_adder_13ccs_18_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_19 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_19_clock),
    .reset(FP_adder_13ccs_19_reset),
    .io_in_a(FP_adder_13ccs_19_io_in_a),
    .io_in_b(FP_adder_13ccs_19_io_in_b),
    .io_out_s(FP_adder_13ccs_19_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_20 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_20_clock),
    .reset(FP_adder_13ccs_20_reset),
    .io_in_a(FP_adder_13ccs_20_io_in_a),
    .io_in_b(FP_adder_13ccs_20_io_in_b),
    .io_out_s(FP_adder_13ccs_20_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_21 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_21_clock),
    .reset(FP_adder_13ccs_21_reset),
    .io_in_a(FP_adder_13ccs_21_io_in_a),
    .io_in_b(FP_adder_13ccs_21_io_in_b),
    .io_out_s(FP_adder_13ccs_21_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_22 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_22_clock),
    .reset(FP_adder_13ccs_22_reset),
    .io_in_a(FP_adder_13ccs_22_io_in_a),
    .io_in_b(FP_adder_13ccs_22_io_in_b),
    .io_out_s(FP_adder_13ccs_22_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_23 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_23_clock),
    .reset(FP_adder_13ccs_23_reset),
    .io_in_a(FP_adder_13ccs_23_io_in_a),
    .io_in_b(FP_adder_13ccs_23_io_in_b),
    .io_out_s(FP_adder_13ccs_23_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_24 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_24_clock),
    .reset(FP_adder_13ccs_24_reset),
    .io_in_a(FP_adder_13ccs_24_io_in_a),
    .io_in_b(FP_adder_13ccs_24_io_in_b),
    .io_out_s(FP_adder_13ccs_24_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_25 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_25_clock),
    .reset(FP_adder_13ccs_25_reset),
    .io_in_a(FP_adder_13ccs_25_io_in_a),
    .io_in_b(FP_adder_13ccs_25_io_in_b),
    .io_out_s(FP_adder_13ccs_25_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_26 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_26_clock),
    .reset(FP_adder_13ccs_26_reset),
    .io_in_a(FP_adder_13ccs_26_io_in_a),
    .io_in_b(FP_adder_13ccs_26_io_in_b),
    .io_out_s(FP_adder_13ccs_26_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_27 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_27_clock),
    .reset(FP_adder_13ccs_27_reset),
    .io_in_a(FP_adder_13ccs_27_io_in_a),
    .io_in_b(FP_adder_13ccs_27_io_in_b),
    .io_out_s(FP_adder_13ccs_27_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_28 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_28_clock),
    .reset(FP_adder_13ccs_28_reset),
    .io_in_a(FP_adder_13ccs_28_io_in_a),
    .io_in_b(FP_adder_13ccs_28_io_in_b),
    .io_out_s(FP_adder_13ccs_28_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_29 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_29_clock),
    .reset(FP_adder_13ccs_29_reset),
    .io_in_a(FP_adder_13ccs_29_io_in_a),
    .io_in_b(FP_adder_13ccs_29_io_in_b),
    .io_out_s(FP_adder_13ccs_29_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_30 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_30_clock),
    .reset(FP_adder_13ccs_30_reset),
    .io_in_a(FP_adder_13ccs_30_io_in_a),
    .io_in_b(FP_adder_13ccs_30_io_in_b),
    .io_out_s(FP_adder_13ccs_30_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_31 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_31_clock),
    .reset(FP_adder_13ccs_31_reset),
    .io_in_a(FP_adder_13ccs_31_io_in_a),
    .io_in_b(FP_adder_13ccs_31_io_in_b),
    .io_out_s(FP_adder_13ccs_31_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_32 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_32_clock),
    .reset(FP_adder_13ccs_32_reset),
    .io_in_a(FP_adder_13ccs_32_io_in_a),
    .io_in_b(FP_adder_13ccs_32_io_in_b),
    .io_out_s(FP_adder_13ccs_32_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_33 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_33_clock),
    .reset(FP_adder_13ccs_33_reset),
    .io_in_a(FP_adder_13ccs_33_io_in_a),
    .io_in_b(FP_adder_13ccs_33_io_in_b),
    .io_out_s(FP_adder_13ccs_33_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_34 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_34_clock),
    .reset(FP_adder_13ccs_34_reset),
    .io_in_a(FP_adder_13ccs_34_io_in_a),
    .io_in_b(FP_adder_13ccs_34_io_in_b),
    .io_out_s(FP_adder_13ccs_34_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_35 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_35_clock),
    .reset(FP_adder_13ccs_35_reset),
    .io_in_a(FP_adder_13ccs_35_io_in_a),
    .io_in_b(FP_adder_13ccs_35_io_in_b),
    .io_out_s(FP_adder_13ccs_35_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_36 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_36_clock),
    .reset(FP_adder_13ccs_36_reset),
    .io_in_a(FP_adder_13ccs_36_io_in_a),
    .io_in_b(FP_adder_13ccs_36_io_in_b),
    .io_out_s(FP_adder_13ccs_36_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_37 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_37_clock),
    .reset(FP_adder_13ccs_37_reset),
    .io_in_a(FP_adder_13ccs_37_io_in_a),
    .io_in_b(FP_adder_13ccs_37_io_in_b),
    .io_out_s(FP_adder_13ccs_37_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_38 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_38_clock),
    .reset(FP_adder_13ccs_38_reset),
    .io_in_a(FP_adder_13ccs_38_io_in_a),
    .io_in_b(FP_adder_13ccs_38_io_in_b),
    .io_out_s(FP_adder_13ccs_38_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_39 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_39_clock),
    .reset(FP_adder_13ccs_39_reset),
    .io_in_a(FP_adder_13ccs_39_io_in_a),
    .io_in_b(FP_adder_13ccs_39_io_in_b),
    .io_out_s(FP_adder_13ccs_39_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_40 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_40_clock),
    .reset(FP_adder_13ccs_40_reset),
    .io_in_a(FP_adder_13ccs_40_io_in_a),
    .io_in_b(FP_adder_13ccs_40_io_in_b),
    .io_out_s(FP_adder_13ccs_40_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_41 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_41_clock),
    .reset(FP_adder_13ccs_41_reset),
    .io_in_a(FP_adder_13ccs_41_io_in_a),
    .io_in_b(FP_adder_13ccs_41_io_in_b),
    .io_out_s(FP_adder_13ccs_41_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_42 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_42_clock),
    .reset(FP_adder_13ccs_42_reset),
    .io_in_a(FP_adder_13ccs_42_io_in_a),
    .io_in_b(FP_adder_13ccs_42_io_in_b),
    .io_out_s(FP_adder_13ccs_42_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_43 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_43_clock),
    .reset(FP_adder_13ccs_43_reset),
    .io_in_a(FP_adder_13ccs_43_io_in_a),
    .io_in_b(FP_adder_13ccs_43_io_in_b),
    .io_out_s(FP_adder_13ccs_43_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_44 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_44_clock),
    .reset(FP_adder_13ccs_44_reset),
    .io_in_a(FP_adder_13ccs_44_io_in_a),
    .io_in_b(FP_adder_13ccs_44_io_in_b),
    .io_out_s(FP_adder_13ccs_44_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_45 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_45_clock),
    .reset(FP_adder_13ccs_45_reset),
    .io_in_a(FP_adder_13ccs_45_io_in_a),
    .io_in_b(FP_adder_13ccs_45_io_in_b),
    .io_out_s(FP_adder_13ccs_45_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_46 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_46_clock),
    .reset(FP_adder_13ccs_46_reset),
    .io_in_a(FP_adder_13ccs_46_io_in_a),
    .io_in_b(FP_adder_13ccs_46_io_in_b),
    .io_out_s(FP_adder_13ccs_46_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_47 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_47_clock),
    .reset(FP_adder_13ccs_47_reset),
    .io_in_a(FP_adder_13ccs_47_io_in_a),
    .io_in_b(FP_adder_13ccs_47_io_in_b),
    .io_out_s(FP_adder_13ccs_47_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_48 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_48_clock),
    .reset(FP_adder_13ccs_48_reset),
    .io_in_a(FP_adder_13ccs_48_io_in_a),
    .io_in_b(FP_adder_13ccs_48_io_in_b),
    .io_out_s(FP_adder_13ccs_48_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_49 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_49_clock),
    .reset(FP_adder_13ccs_49_reset),
    .io_in_a(FP_adder_13ccs_49_io_in_a),
    .io_in_b(FP_adder_13ccs_49_io_in_b),
    .io_out_s(FP_adder_13ccs_49_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_50 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_50_clock),
    .reset(FP_adder_13ccs_50_reset),
    .io_in_a(FP_adder_13ccs_50_io_in_a),
    .io_in_b(FP_adder_13ccs_50_io_in_b),
    .io_out_s(FP_adder_13ccs_50_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_51 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_51_clock),
    .reset(FP_adder_13ccs_51_reset),
    .io_in_a(FP_adder_13ccs_51_io_in_a),
    .io_in_b(FP_adder_13ccs_51_io_in_b),
    .io_out_s(FP_adder_13ccs_51_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_52 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_52_clock),
    .reset(FP_adder_13ccs_52_reset),
    .io_in_a(FP_adder_13ccs_52_io_in_a),
    .io_in_b(FP_adder_13ccs_52_io_in_b),
    .io_out_s(FP_adder_13ccs_52_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_53 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_53_clock),
    .reset(FP_adder_13ccs_53_reset),
    .io_in_a(FP_adder_13ccs_53_io_in_a),
    .io_in_b(FP_adder_13ccs_53_io_in_b),
    .io_out_s(FP_adder_13ccs_53_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_54 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_54_clock),
    .reset(FP_adder_13ccs_54_reset),
    .io_in_a(FP_adder_13ccs_54_io_in_a),
    .io_in_b(FP_adder_13ccs_54_io_in_b),
    .io_out_s(FP_adder_13ccs_54_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_55 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_55_clock),
    .reset(FP_adder_13ccs_55_reset),
    .io_in_a(FP_adder_13ccs_55_io_in_a),
    .io_in_b(FP_adder_13ccs_55_io_in_b),
    .io_out_s(FP_adder_13ccs_55_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_56 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_56_clock),
    .reset(FP_adder_13ccs_56_reset),
    .io_in_a(FP_adder_13ccs_56_io_in_a),
    .io_in_b(FP_adder_13ccs_56_io_in_b),
    .io_out_s(FP_adder_13ccs_56_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_57 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_57_clock),
    .reset(FP_adder_13ccs_57_reset),
    .io_in_a(FP_adder_13ccs_57_io_in_a),
    .io_in_b(FP_adder_13ccs_57_io_in_b),
    .io_out_s(FP_adder_13ccs_57_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_58 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_58_clock),
    .reset(FP_adder_13ccs_58_reset),
    .io_in_a(FP_adder_13ccs_58_io_in_a),
    .io_in_b(FP_adder_13ccs_58_io_in_b),
    .io_out_s(FP_adder_13ccs_58_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_59 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_59_clock),
    .reset(FP_adder_13ccs_59_reset),
    .io_in_a(FP_adder_13ccs_59_io_in_a),
    .io_in_b(FP_adder_13ccs_59_io_in_b),
    .io_out_s(FP_adder_13ccs_59_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_60 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_60_clock),
    .reset(FP_adder_13ccs_60_reset),
    .io_in_a(FP_adder_13ccs_60_io_in_a),
    .io_in_b(FP_adder_13ccs_60_io_in_b),
    .io_out_s(FP_adder_13ccs_60_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_61 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_61_clock),
    .reset(FP_adder_13ccs_61_reset),
    .io_in_a(FP_adder_13ccs_61_io_in_a),
    .io_in_b(FP_adder_13ccs_61_io_in_b),
    .io_out_s(FP_adder_13ccs_61_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_62 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_62_clock),
    .reset(FP_adder_13ccs_62_reset),
    .io_in_a(FP_adder_13ccs_62_io_in_a),
    .io_in_b(FP_adder_13ccs_62_io_in_b),
    .io_out_s(FP_adder_13ccs_62_io_out_s)
  );
  FP_adder_13ccs FP_adder_13ccs_63 ( // @[FloatingPointDesigns.scala 2490:25]
    .clock(FP_adder_13ccs_63_clock),
    .reset(FP_adder_13ccs_63_reset),
    .io_in_a(FP_adder_13ccs_63_io_in_a),
    .io_in_b(FP_adder_13ccs_63_io_in_b),
    .io_out_s(FP_adder_13ccs_63_io_out_s)
  );
  FPReg FPReg ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_clock),
    .reset(FPReg_reset),
    .io_in(FPReg_io_in),
    .io_out(FPReg_io_out)
  );
  FPReg FPReg_1 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_1_clock),
    .reset(FPReg_1_reset),
    .io_in(FPReg_1_io_in),
    .io_out(FPReg_1_io_out)
  );
  FPReg FPReg_2 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_2_clock),
    .reset(FPReg_2_reset),
    .io_in(FPReg_2_io_in),
    .io_out(FPReg_2_io_out)
  );
  FPReg FPReg_3 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_3_clock),
    .reset(FPReg_3_reset),
    .io_in(FPReg_3_io_in),
    .io_out(FPReg_3_io_out)
  );
  FPReg FPReg_4 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_4_clock),
    .reset(FPReg_4_reset),
    .io_in(FPReg_4_io_in),
    .io_out(FPReg_4_io_out)
  );
  FPReg FPReg_5 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_5_clock),
    .reset(FPReg_5_reset),
    .io_in(FPReg_5_io_in),
    .io_out(FPReg_5_io_out)
  );
  FPReg FPReg_6 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_6_clock),
    .reset(FPReg_6_reset),
    .io_in(FPReg_6_io_in),
    .io_out(FPReg_6_io_out)
  );
  FPReg FPReg_7 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_7_clock),
    .reset(FPReg_7_reset),
    .io_in(FPReg_7_io_in),
    .io_out(FPReg_7_io_out)
  );
  FPReg FPReg_8 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_8_clock),
    .reset(FPReg_8_reset),
    .io_in(FPReg_8_io_in),
    .io_out(FPReg_8_io_out)
  );
  FPReg FPReg_9 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_9_clock),
    .reset(FPReg_9_reset),
    .io_in(FPReg_9_io_in),
    .io_out(FPReg_9_io_out)
  );
  FPReg FPReg_10 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_10_clock),
    .reset(FPReg_10_reset),
    .io_in(FPReg_10_io_in),
    .io_out(FPReg_10_io_out)
  );
  FPReg FPReg_11 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_11_clock),
    .reset(FPReg_11_reset),
    .io_in(FPReg_11_io_in),
    .io_out(FPReg_11_io_out)
  );
  FPReg FPReg_12 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_12_clock),
    .reset(FPReg_12_reset),
    .io_in(FPReg_12_io_in),
    .io_out(FPReg_12_io_out)
  );
  FPReg FPReg_13 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_13_clock),
    .reset(FPReg_13_reset),
    .io_in(FPReg_13_io_in),
    .io_out(FPReg_13_io_out)
  );
  FPReg FPReg_14 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_14_clock),
    .reset(FPReg_14_reset),
    .io_in(FPReg_14_io_in),
    .io_out(FPReg_14_io_out)
  );
  FPReg FPReg_15 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_15_clock),
    .reset(FPReg_15_reset),
    .io_in(FPReg_15_io_in),
    .io_out(FPReg_15_io_out)
  );
  FPReg FPReg_16 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_16_clock),
    .reset(FPReg_16_reset),
    .io_in(FPReg_16_io_in),
    .io_out(FPReg_16_io_out)
  );
  FPReg FPReg_17 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_17_clock),
    .reset(FPReg_17_reset),
    .io_in(FPReg_17_io_in),
    .io_out(FPReg_17_io_out)
  );
  FPReg FPReg_18 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_18_clock),
    .reset(FPReg_18_reset),
    .io_in(FPReg_18_io_in),
    .io_out(FPReg_18_io_out)
  );
  FPReg FPReg_19 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_19_clock),
    .reset(FPReg_19_reset),
    .io_in(FPReg_19_io_in),
    .io_out(FPReg_19_io_out)
  );
  FPReg FPReg_20 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_20_clock),
    .reset(FPReg_20_reset),
    .io_in(FPReg_20_io_in),
    .io_out(FPReg_20_io_out)
  );
  FPReg FPReg_21 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_21_clock),
    .reset(FPReg_21_reset),
    .io_in(FPReg_21_io_in),
    .io_out(FPReg_21_io_out)
  );
  FPReg FPReg_22 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_22_clock),
    .reset(FPReg_22_reset),
    .io_in(FPReg_22_io_in),
    .io_out(FPReg_22_io_out)
  );
  FPReg FPReg_23 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_23_clock),
    .reset(FPReg_23_reset),
    .io_in(FPReg_23_io_in),
    .io_out(FPReg_23_io_out)
  );
  FPReg FPReg_24 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_24_clock),
    .reset(FPReg_24_reset),
    .io_in(FPReg_24_io_in),
    .io_out(FPReg_24_io_out)
  );
  FPReg FPReg_25 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_25_clock),
    .reset(FPReg_25_reset),
    .io_in(FPReg_25_io_in),
    .io_out(FPReg_25_io_out)
  );
  FPReg FPReg_26 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_26_clock),
    .reset(FPReg_26_reset),
    .io_in(FPReg_26_io_in),
    .io_out(FPReg_26_io_out)
  );
  FPReg FPReg_27 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_27_clock),
    .reset(FPReg_27_reset),
    .io_in(FPReg_27_io_in),
    .io_out(FPReg_27_io_out)
  );
  FPReg FPReg_28 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_28_clock),
    .reset(FPReg_28_reset),
    .io_in(FPReg_28_io_in),
    .io_out(FPReg_28_io_out)
  );
  FPReg FPReg_29 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_29_clock),
    .reset(FPReg_29_reset),
    .io_in(FPReg_29_io_in),
    .io_out(FPReg_29_io_out)
  );
  FPReg FPReg_30 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_30_clock),
    .reset(FPReg_30_reset),
    .io_in(FPReg_30_io_in),
    .io_out(FPReg_30_io_out)
  );
  FPReg FPReg_31 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_31_clock),
    .reset(FPReg_31_reset),
    .io_in(FPReg_31_io_in),
    .io_out(FPReg_31_io_out)
  );
  FPReg FPReg_32 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_32_clock),
    .reset(FPReg_32_reset),
    .io_in(FPReg_32_io_in),
    .io_out(FPReg_32_io_out)
  );
  FPReg FPReg_33 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_33_clock),
    .reset(FPReg_33_reset),
    .io_in(FPReg_33_io_in),
    .io_out(FPReg_33_io_out)
  );
  FPReg FPReg_34 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_34_clock),
    .reset(FPReg_34_reset),
    .io_in(FPReg_34_io_in),
    .io_out(FPReg_34_io_out)
  );
  FPReg FPReg_35 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_35_clock),
    .reset(FPReg_35_reset),
    .io_in(FPReg_35_io_in),
    .io_out(FPReg_35_io_out)
  );
  FPReg FPReg_36 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_36_clock),
    .reset(FPReg_36_reset),
    .io_in(FPReg_36_io_in),
    .io_out(FPReg_36_io_out)
  );
  FPReg FPReg_37 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_37_clock),
    .reset(FPReg_37_reset),
    .io_in(FPReg_37_io_in),
    .io_out(FPReg_37_io_out)
  );
  FPReg FPReg_38 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_38_clock),
    .reset(FPReg_38_reset),
    .io_in(FPReg_38_io_in),
    .io_out(FPReg_38_io_out)
  );
  FPReg FPReg_39 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_39_clock),
    .reset(FPReg_39_reset),
    .io_in(FPReg_39_io_in),
    .io_out(FPReg_39_io_out)
  );
  FPReg FPReg_40 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_40_clock),
    .reset(FPReg_40_reset),
    .io_in(FPReg_40_io_in),
    .io_out(FPReg_40_io_out)
  );
  FPReg FPReg_41 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_41_clock),
    .reset(FPReg_41_reset),
    .io_in(FPReg_41_io_in),
    .io_out(FPReg_41_io_out)
  );
  FPReg FPReg_42 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_42_clock),
    .reset(FPReg_42_reset),
    .io_in(FPReg_42_io_in),
    .io_out(FPReg_42_io_out)
  );
  FPReg FPReg_43 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_43_clock),
    .reset(FPReg_43_reset),
    .io_in(FPReg_43_io_in),
    .io_out(FPReg_43_io_out)
  );
  FPReg FPReg_44 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_44_clock),
    .reset(FPReg_44_reset),
    .io_in(FPReg_44_io_in),
    .io_out(FPReg_44_io_out)
  );
  FPReg FPReg_45 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_45_clock),
    .reset(FPReg_45_reset),
    .io_in(FPReg_45_io_in),
    .io_out(FPReg_45_io_out)
  );
  FPReg FPReg_46 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_46_clock),
    .reset(FPReg_46_reset),
    .io_in(FPReg_46_io_in),
    .io_out(FPReg_46_io_out)
  );
  FPReg FPReg_47 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_47_clock),
    .reset(FPReg_47_reset),
    .io_in(FPReg_47_io_in),
    .io_out(FPReg_47_io_out)
  );
  FPReg FPReg_48 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_48_clock),
    .reset(FPReg_48_reset),
    .io_in(FPReg_48_io_in),
    .io_out(FPReg_48_io_out)
  );
  FPReg FPReg_49 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_49_clock),
    .reset(FPReg_49_reset),
    .io_in(FPReg_49_io_in),
    .io_out(FPReg_49_io_out)
  );
  FPReg FPReg_50 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_50_clock),
    .reset(FPReg_50_reset),
    .io_in(FPReg_50_io_in),
    .io_out(FPReg_50_io_out)
  );
  FPReg FPReg_51 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_51_clock),
    .reset(FPReg_51_reset),
    .io_in(FPReg_51_io_in),
    .io_out(FPReg_51_io_out)
  );
  FPReg FPReg_52 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_52_clock),
    .reset(FPReg_52_reset),
    .io_in(FPReg_52_io_in),
    .io_out(FPReg_52_io_out)
  );
  FPReg FPReg_53 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_53_clock),
    .reset(FPReg_53_reset),
    .io_in(FPReg_53_io_in),
    .io_out(FPReg_53_io_out)
  );
  FPReg FPReg_54 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_54_clock),
    .reset(FPReg_54_reset),
    .io_in(FPReg_54_io_in),
    .io_out(FPReg_54_io_out)
  );
  FPReg FPReg_55 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_55_clock),
    .reset(FPReg_55_reset),
    .io_in(FPReg_55_io_in),
    .io_out(FPReg_55_io_out)
  );
  FPReg FPReg_56 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_56_clock),
    .reset(FPReg_56_reset),
    .io_in(FPReg_56_io_in),
    .io_out(FPReg_56_io_out)
  );
  FPReg FPReg_57 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_57_clock),
    .reset(FPReg_57_reset),
    .io_in(FPReg_57_io_in),
    .io_out(FPReg_57_io_out)
  );
  FPReg FPReg_58 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_58_clock),
    .reset(FPReg_58_reset),
    .io_in(FPReg_58_io_in),
    .io_out(FPReg_58_io_out)
  );
  FPReg FPReg_59 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_59_clock),
    .reset(FPReg_59_reset),
    .io_in(FPReg_59_io_in),
    .io_out(FPReg_59_io_out)
  );
  FPReg FPReg_60 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_60_clock),
    .reset(FPReg_60_reset),
    .io_in(FPReg_60_io_in),
    .io_out(FPReg_60_io_out)
  );
  FPReg FPReg_61 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_61_clock),
    .reset(FPReg_61_reset),
    .io_in(FPReg_61_io_in),
    .io_out(FPReg_61_io_out)
  );
  FPReg FPReg_62 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_62_clock),
    .reset(FPReg_62_reset),
    .io_in(FPReg_62_io_in),
    .io_out(FPReg_62_io_out)
  );
  FPReg FPReg_63 ( // @[FloatingPointDesigns.scala 2494:48]
    .clock(FPReg_63_clock),
    .reset(FPReg_63_reset),
    .io_in(FPReg_63_io_in),
    .io_out(FPReg_63_io_out)
  );
  assign io_out_s_0 = FP_adder_13ccs_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_1 = FP_adder_13ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_2 = FP_adder_13ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_3 = FP_adder_13ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_4 = FP_adder_13ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_5 = FP_adder_13ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_6 = FP_adder_13ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_7 = FP_adder_13ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_8 = FP_adder_13ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_9 = FP_adder_13ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_10 = FP_adder_13ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_11 = FP_adder_13ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_12 = FP_adder_13ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_13 = FP_adder_13ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_14 = FP_adder_13ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_15 = FP_adder_13ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_16 = FP_adder_13ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_17 = FP_adder_13ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_18 = FP_adder_13ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_19 = FP_adder_13ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_20 = FP_adder_13ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_21 = FP_adder_13ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_22 = FP_adder_13ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_23 = FP_adder_13ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_24 = FP_adder_13ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_25 = FP_adder_13ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_26 = FP_adder_13ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_27 = FP_adder_13ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_28 = FP_adder_13ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_29 = FP_adder_13ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_30 = FP_adder_13ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_31 = FP_adder_13ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_32 = FP_adder_13ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_33 = FP_adder_13ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_34 = FP_adder_13ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_35 = FP_adder_13ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_36 = FP_adder_13ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_37 = FP_adder_13ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_38 = FP_adder_13ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_39 = FP_adder_13ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_40 = FP_adder_13ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_41 = FP_adder_13ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_42 = FP_adder_13ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_43 = FP_adder_13ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_44 = FP_adder_13ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_45 = FP_adder_13ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_46 = FP_adder_13ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_47 = FP_adder_13ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_48 = FP_adder_13ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_49 = FP_adder_13ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_50 = FP_adder_13ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_51 = FP_adder_13ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_52 = FP_adder_13ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_53 = FP_adder_13ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_54 = FP_adder_13ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_55 = FP_adder_13ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_56 = FP_adder_13ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_57 = FP_adder_13ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_58 = FP_adder_13ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_59 = FP_adder_13ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_60 = FP_adder_13ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_61 = FP_adder_13ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_62 = FP_adder_13ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign io_out_s_63 = FP_adder_13ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2501:19]
  assign FP_multiplier_10ccs_clock = clock;
  assign FP_multiplier_10ccs_reset = reset;
  assign FP_multiplier_10ccs_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_io_in_b = io_in_b_0; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_1_clock = clock;
  assign FP_multiplier_10ccs_1_reset = reset;
  assign FP_multiplier_10ccs_1_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_1_io_in_b = io_in_b_1; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_2_clock = clock;
  assign FP_multiplier_10ccs_2_reset = reset;
  assign FP_multiplier_10ccs_2_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_2_io_in_b = io_in_b_2; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_3_clock = clock;
  assign FP_multiplier_10ccs_3_reset = reset;
  assign FP_multiplier_10ccs_3_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_3_io_in_b = io_in_b_3; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_4_clock = clock;
  assign FP_multiplier_10ccs_4_reset = reset;
  assign FP_multiplier_10ccs_4_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_4_io_in_b = io_in_b_4; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_5_clock = clock;
  assign FP_multiplier_10ccs_5_reset = reset;
  assign FP_multiplier_10ccs_5_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_5_io_in_b = io_in_b_5; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_6_clock = clock;
  assign FP_multiplier_10ccs_6_reset = reset;
  assign FP_multiplier_10ccs_6_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_6_io_in_b = io_in_b_6; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_7_clock = clock;
  assign FP_multiplier_10ccs_7_reset = reset;
  assign FP_multiplier_10ccs_7_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_7_io_in_b = io_in_b_7; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_8_clock = clock;
  assign FP_multiplier_10ccs_8_reset = reset;
  assign FP_multiplier_10ccs_8_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_8_io_in_b = io_in_b_8; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_9_clock = clock;
  assign FP_multiplier_10ccs_9_reset = reset;
  assign FP_multiplier_10ccs_9_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_9_io_in_b = io_in_b_9; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_10_clock = clock;
  assign FP_multiplier_10ccs_10_reset = reset;
  assign FP_multiplier_10ccs_10_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_10_io_in_b = io_in_b_10; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_11_clock = clock;
  assign FP_multiplier_10ccs_11_reset = reset;
  assign FP_multiplier_10ccs_11_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_11_io_in_b = io_in_b_11; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_12_clock = clock;
  assign FP_multiplier_10ccs_12_reset = reset;
  assign FP_multiplier_10ccs_12_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_12_io_in_b = io_in_b_12; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_13_clock = clock;
  assign FP_multiplier_10ccs_13_reset = reset;
  assign FP_multiplier_10ccs_13_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_13_io_in_b = io_in_b_13; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_14_clock = clock;
  assign FP_multiplier_10ccs_14_reset = reset;
  assign FP_multiplier_10ccs_14_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_14_io_in_b = io_in_b_14; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_15_clock = clock;
  assign FP_multiplier_10ccs_15_reset = reset;
  assign FP_multiplier_10ccs_15_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_15_io_in_b = io_in_b_15; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_16_clock = clock;
  assign FP_multiplier_10ccs_16_reset = reset;
  assign FP_multiplier_10ccs_16_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_16_io_in_b = io_in_b_16; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_17_clock = clock;
  assign FP_multiplier_10ccs_17_reset = reset;
  assign FP_multiplier_10ccs_17_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_17_io_in_b = io_in_b_17; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_18_clock = clock;
  assign FP_multiplier_10ccs_18_reset = reset;
  assign FP_multiplier_10ccs_18_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_18_io_in_b = io_in_b_18; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_19_clock = clock;
  assign FP_multiplier_10ccs_19_reset = reset;
  assign FP_multiplier_10ccs_19_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_19_io_in_b = io_in_b_19; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_20_clock = clock;
  assign FP_multiplier_10ccs_20_reset = reset;
  assign FP_multiplier_10ccs_20_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_20_io_in_b = io_in_b_20; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_21_clock = clock;
  assign FP_multiplier_10ccs_21_reset = reset;
  assign FP_multiplier_10ccs_21_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_21_io_in_b = io_in_b_21; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_22_clock = clock;
  assign FP_multiplier_10ccs_22_reset = reset;
  assign FP_multiplier_10ccs_22_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_22_io_in_b = io_in_b_22; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_23_clock = clock;
  assign FP_multiplier_10ccs_23_reset = reset;
  assign FP_multiplier_10ccs_23_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_23_io_in_b = io_in_b_23; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_24_clock = clock;
  assign FP_multiplier_10ccs_24_reset = reset;
  assign FP_multiplier_10ccs_24_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_24_io_in_b = io_in_b_24; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_25_clock = clock;
  assign FP_multiplier_10ccs_25_reset = reset;
  assign FP_multiplier_10ccs_25_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_25_io_in_b = io_in_b_25; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_26_clock = clock;
  assign FP_multiplier_10ccs_26_reset = reset;
  assign FP_multiplier_10ccs_26_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_26_io_in_b = io_in_b_26; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_27_clock = clock;
  assign FP_multiplier_10ccs_27_reset = reset;
  assign FP_multiplier_10ccs_27_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_27_io_in_b = io_in_b_27; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_28_clock = clock;
  assign FP_multiplier_10ccs_28_reset = reset;
  assign FP_multiplier_10ccs_28_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_28_io_in_b = io_in_b_28; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_29_clock = clock;
  assign FP_multiplier_10ccs_29_reset = reset;
  assign FP_multiplier_10ccs_29_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_29_io_in_b = io_in_b_29; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_30_clock = clock;
  assign FP_multiplier_10ccs_30_reset = reset;
  assign FP_multiplier_10ccs_30_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_30_io_in_b = io_in_b_30; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_31_clock = clock;
  assign FP_multiplier_10ccs_31_reset = reset;
  assign FP_multiplier_10ccs_31_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_31_io_in_b = io_in_b_31; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_32_clock = clock;
  assign FP_multiplier_10ccs_32_reset = reset;
  assign FP_multiplier_10ccs_32_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_32_io_in_b = io_in_b_32; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_33_clock = clock;
  assign FP_multiplier_10ccs_33_reset = reset;
  assign FP_multiplier_10ccs_33_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_33_io_in_b = io_in_b_33; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_34_clock = clock;
  assign FP_multiplier_10ccs_34_reset = reset;
  assign FP_multiplier_10ccs_34_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_34_io_in_b = io_in_b_34; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_35_clock = clock;
  assign FP_multiplier_10ccs_35_reset = reset;
  assign FP_multiplier_10ccs_35_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_35_io_in_b = io_in_b_35; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_36_clock = clock;
  assign FP_multiplier_10ccs_36_reset = reset;
  assign FP_multiplier_10ccs_36_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_36_io_in_b = io_in_b_36; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_37_clock = clock;
  assign FP_multiplier_10ccs_37_reset = reset;
  assign FP_multiplier_10ccs_37_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_37_io_in_b = io_in_b_37; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_38_clock = clock;
  assign FP_multiplier_10ccs_38_reset = reset;
  assign FP_multiplier_10ccs_38_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_38_io_in_b = io_in_b_38; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_39_clock = clock;
  assign FP_multiplier_10ccs_39_reset = reset;
  assign FP_multiplier_10ccs_39_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_39_io_in_b = io_in_b_39; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_40_clock = clock;
  assign FP_multiplier_10ccs_40_reset = reset;
  assign FP_multiplier_10ccs_40_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_40_io_in_b = io_in_b_40; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_41_clock = clock;
  assign FP_multiplier_10ccs_41_reset = reset;
  assign FP_multiplier_10ccs_41_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_41_io_in_b = io_in_b_41; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_42_clock = clock;
  assign FP_multiplier_10ccs_42_reset = reset;
  assign FP_multiplier_10ccs_42_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_42_io_in_b = io_in_b_42; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_43_clock = clock;
  assign FP_multiplier_10ccs_43_reset = reset;
  assign FP_multiplier_10ccs_43_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_43_io_in_b = io_in_b_43; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_44_clock = clock;
  assign FP_multiplier_10ccs_44_reset = reset;
  assign FP_multiplier_10ccs_44_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_44_io_in_b = io_in_b_44; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_45_clock = clock;
  assign FP_multiplier_10ccs_45_reset = reset;
  assign FP_multiplier_10ccs_45_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_45_io_in_b = io_in_b_45; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_46_clock = clock;
  assign FP_multiplier_10ccs_46_reset = reset;
  assign FP_multiplier_10ccs_46_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_46_io_in_b = io_in_b_46; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_47_clock = clock;
  assign FP_multiplier_10ccs_47_reset = reset;
  assign FP_multiplier_10ccs_47_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_47_io_in_b = io_in_b_47; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_48_clock = clock;
  assign FP_multiplier_10ccs_48_reset = reset;
  assign FP_multiplier_10ccs_48_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_48_io_in_b = io_in_b_48; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_49_clock = clock;
  assign FP_multiplier_10ccs_49_reset = reset;
  assign FP_multiplier_10ccs_49_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_49_io_in_b = io_in_b_49; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_50_clock = clock;
  assign FP_multiplier_10ccs_50_reset = reset;
  assign FP_multiplier_10ccs_50_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_50_io_in_b = io_in_b_50; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_51_clock = clock;
  assign FP_multiplier_10ccs_51_reset = reset;
  assign FP_multiplier_10ccs_51_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_51_io_in_b = io_in_b_51; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_52_clock = clock;
  assign FP_multiplier_10ccs_52_reset = reset;
  assign FP_multiplier_10ccs_52_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_52_io_in_b = io_in_b_52; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_53_clock = clock;
  assign FP_multiplier_10ccs_53_reset = reset;
  assign FP_multiplier_10ccs_53_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_53_io_in_b = io_in_b_53; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_54_clock = clock;
  assign FP_multiplier_10ccs_54_reset = reset;
  assign FP_multiplier_10ccs_54_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_54_io_in_b = io_in_b_54; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_55_clock = clock;
  assign FP_multiplier_10ccs_55_reset = reset;
  assign FP_multiplier_10ccs_55_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_55_io_in_b = io_in_b_55; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_56_clock = clock;
  assign FP_multiplier_10ccs_56_reset = reset;
  assign FP_multiplier_10ccs_56_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_56_io_in_b = io_in_b_56; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_57_clock = clock;
  assign FP_multiplier_10ccs_57_reset = reset;
  assign FP_multiplier_10ccs_57_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_57_io_in_b = io_in_b_57; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_58_clock = clock;
  assign FP_multiplier_10ccs_58_reset = reset;
  assign FP_multiplier_10ccs_58_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_58_io_in_b = io_in_b_58; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_59_clock = clock;
  assign FP_multiplier_10ccs_59_reset = reset;
  assign FP_multiplier_10ccs_59_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_59_io_in_b = io_in_b_59; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_60_clock = clock;
  assign FP_multiplier_10ccs_60_reset = reset;
  assign FP_multiplier_10ccs_60_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_60_io_in_b = io_in_b_60; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_61_clock = clock;
  assign FP_multiplier_10ccs_61_reset = reset;
  assign FP_multiplier_10ccs_61_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_61_io_in_b = io_in_b_61; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_62_clock = clock;
  assign FP_multiplier_10ccs_62_reset = reset;
  assign FP_multiplier_10ccs_62_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_62_io_in_b = io_in_b_62; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_multiplier_10ccs_63_clock = clock;
  assign FP_multiplier_10ccs_63_reset = reset;
  assign FP_multiplier_10ccs_63_io_in_a = io_in_a; // @[FloatingPointDesigns.scala 2496:30]
  assign FP_multiplier_10ccs_63_io_in_b = io_in_b_63; // @[FloatingPointDesigns.scala 2497:30]
  assign FP_adder_13ccs_clock = clock;
  assign FP_adder_13ccs_reset = reset;
  assign FP_adder_13ccs_io_in_a = FP_multiplier_10ccs_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_io_in_b = FPReg_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_1_clock = clock;
  assign FP_adder_13ccs_1_reset = reset;
  assign FP_adder_13ccs_1_io_in_a = FP_multiplier_10ccs_1_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_1_io_in_b = FPReg_1_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_2_clock = clock;
  assign FP_adder_13ccs_2_reset = reset;
  assign FP_adder_13ccs_2_io_in_a = FP_multiplier_10ccs_2_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_2_io_in_b = FPReg_2_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_3_clock = clock;
  assign FP_adder_13ccs_3_reset = reset;
  assign FP_adder_13ccs_3_io_in_a = FP_multiplier_10ccs_3_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_3_io_in_b = FPReg_3_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_4_clock = clock;
  assign FP_adder_13ccs_4_reset = reset;
  assign FP_adder_13ccs_4_io_in_a = FP_multiplier_10ccs_4_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_4_io_in_b = FPReg_4_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_5_clock = clock;
  assign FP_adder_13ccs_5_reset = reset;
  assign FP_adder_13ccs_5_io_in_a = FP_multiplier_10ccs_5_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_5_io_in_b = FPReg_5_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_6_clock = clock;
  assign FP_adder_13ccs_6_reset = reset;
  assign FP_adder_13ccs_6_io_in_a = FP_multiplier_10ccs_6_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_6_io_in_b = FPReg_6_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_7_clock = clock;
  assign FP_adder_13ccs_7_reset = reset;
  assign FP_adder_13ccs_7_io_in_a = FP_multiplier_10ccs_7_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_7_io_in_b = FPReg_7_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_8_clock = clock;
  assign FP_adder_13ccs_8_reset = reset;
  assign FP_adder_13ccs_8_io_in_a = FP_multiplier_10ccs_8_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_8_io_in_b = FPReg_8_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_9_clock = clock;
  assign FP_adder_13ccs_9_reset = reset;
  assign FP_adder_13ccs_9_io_in_a = FP_multiplier_10ccs_9_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_9_io_in_b = FPReg_9_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_10_clock = clock;
  assign FP_adder_13ccs_10_reset = reset;
  assign FP_adder_13ccs_10_io_in_a = FP_multiplier_10ccs_10_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_10_io_in_b = FPReg_10_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_11_clock = clock;
  assign FP_adder_13ccs_11_reset = reset;
  assign FP_adder_13ccs_11_io_in_a = FP_multiplier_10ccs_11_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_11_io_in_b = FPReg_11_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_12_clock = clock;
  assign FP_adder_13ccs_12_reset = reset;
  assign FP_adder_13ccs_12_io_in_a = FP_multiplier_10ccs_12_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_12_io_in_b = FPReg_12_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_13_clock = clock;
  assign FP_adder_13ccs_13_reset = reset;
  assign FP_adder_13ccs_13_io_in_a = FP_multiplier_10ccs_13_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_13_io_in_b = FPReg_13_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_14_clock = clock;
  assign FP_adder_13ccs_14_reset = reset;
  assign FP_adder_13ccs_14_io_in_a = FP_multiplier_10ccs_14_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_14_io_in_b = FPReg_14_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_15_clock = clock;
  assign FP_adder_13ccs_15_reset = reset;
  assign FP_adder_13ccs_15_io_in_a = FP_multiplier_10ccs_15_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_15_io_in_b = FPReg_15_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_16_clock = clock;
  assign FP_adder_13ccs_16_reset = reset;
  assign FP_adder_13ccs_16_io_in_a = FP_multiplier_10ccs_16_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_16_io_in_b = FPReg_16_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_17_clock = clock;
  assign FP_adder_13ccs_17_reset = reset;
  assign FP_adder_13ccs_17_io_in_a = FP_multiplier_10ccs_17_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_17_io_in_b = FPReg_17_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_18_clock = clock;
  assign FP_adder_13ccs_18_reset = reset;
  assign FP_adder_13ccs_18_io_in_a = FP_multiplier_10ccs_18_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_18_io_in_b = FPReg_18_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_19_clock = clock;
  assign FP_adder_13ccs_19_reset = reset;
  assign FP_adder_13ccs_19_io_in_a = FP_multiplier_10ccs_19_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_19_io_in_b = FPReg_19_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_20_clock = clock;
  assign FP_adder_13ccs_20_reset = reset;
  assign FP_adder_13ccs_20_io_in_a = FP_multiplier_10ccs_20_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_20_io_in_b = FPReg_20_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_21_clock = clock;
  assign FP_adder_13ccs_21_reset = reset;
  assign FP_adder_13ccs_21_io_in_a = FP_multiplier_10ccs_21_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_21_io_in_b = FPReg_21_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_22_clock = clock;
  assign FP_adder_13ccs_22_reset = reset;
  assign FP_adder_13ccs_22_io_in_a = FP_multiplier_10ccs_22_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_22_io_in_b = FPReg_22_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_23_clock = clock;
  assign FP_adder_13ccs_23_reset = reset;
  assign FP_adder_13ccs_23_io_in_a = FP_multiplier_10ccs_23_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_23_io_in_b = FPReg_23_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_24_clock = clock;
  assign FP_adder_13ccs_24_reset = reset;
  assign FP_adder_13ccs_24_io_in_a = FP_multiplier_10ccs_24_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_24_io_in_b = FPReg_24_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_25_clock = clock;
  assign FP_adder_13ccs_25_reset = reset;
  assign FP_adder_13ccs_25_io_in_a = FP_multiplier_10ccs_25_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_25_io_in_b = FPReg_25_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_26_clock = clock;
  assign FP_adder_13ccs_26_reset = reset;
  assign FP_adder_13ccs_26_io_in_a = FP_multiplier_10ccs_26_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_26_io_in_b = FPReg_26_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_27_clock = clock;
  assign FP_adder_13ccs_27_reset = reset;
  assign FP_adder_13ccs_27_io_in_a = FP_multiplier_10ccs_27_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_27_io_in_b = FPReg_27_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_28_clock = clock;
  assign FP_adder_13ccs_28_reset = reset;
  assign FP_adder_13ccs_28_io_in_a = FP_multiplier_10ccs_28_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_28_io_in_b = FPReg_28_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_29_clock = clock;
  assign FP_adder_13ccs_29_reset = reset;
  assign FP_adder_13ccs_29_io_in_a = FP_multiplier_10ccs_29_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_29_io_in_b = FPReg_29_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_30_clock = clock;
  assign FP_adder_13ccs_30_reset = reset;
  assign FP_adder_13ccs_30_io_in_a = FP_multiplier_10ccs_30_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_30_io_in_b = FPReg_30_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_31_clock = clock;
  assign FP_adder_13ccs_31_reset = reset;
  assign FP_adder_13ccs_31_io_in_a = FP_multiplier_10ccs_31_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_31_io_in_b = FPReg_31_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_32_clock = clock;
  assign FP_adder_13ccs_32_reset = reset;
  assign FP_adder_13ccs_32_io_in_a = FP_multiplier_10ccs_32_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_32_io_in_b = FPReg_32_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_33_clock = clock;
  assign FP_adder_13ccs_33_reset = reset;
  assign FP_adder_13ccs_33_io_in_a = FP_multiplier_10ccs_33_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_33_io_in_b = FPReg_33_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_34_clock = clock;
  assign FP_adder_13ccs_34_reset = reset;
  assign FP_adder_13ccs_34_io_in_a = FP_multiplier_10ccs_34_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_34_io_in_b = FPReg_34_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_35_clock = clock;
  assign FP_adder_13ccs_35_reset = reset;
  assign FP_adder_13ccs_35_io_in_a = FP_multiplier_10ccs_35_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_35_io_in_b = FPReg_35_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_36_clock = clock;
  assign FP_adder_13ccs_36_reset = reset;
  assign FP_adder_13ccs_36_io_in_a = FP_multiplier_10ccs_36_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_36_io_in_b = FPReg_36_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_37_clock = clock;
  assign FP_adder_13ccs_37_reset = reset;
  assign FP_adder_13ccs_37_io_in_a = FP_multiplier_10ccs_37_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_37_io_in_b = FPReg_37_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_38_clock = clock;
  assign FP_adder_13ccs_38_reset = reset;
  assign FP_adder_13ccs_38_io_in_a = FP_multiplier_10ccs_38_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_38_io_in_b = FPReg_38_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_39_clock = clock;
  assign FP_adder_13ccs_39_reset = reset;
  assign FP_adder_13ccs_39_io_in_a = FP_multiplier_10ccs_39_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_39_io_in_b = FPReg_39_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_40_clock = clock;
  assign FP_adder_13ccs_40_reset = reset;
  assign FP_adder_13ccs_40_io_in_a = FP_multiplier_10ccs_40_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_40_io_in_b = FPReg_40_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_41_clock = clock;
  assign FP_adder_13ccs_41_reset = reset;
  assign FP_adder_13ccs_41_io_in_a = FP_multiplier_10ccs_41_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_41_io_in_b = FPReg_41_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_42_clock = clock;
  assign FP_adder_13ccs_42_reset = reset;
  assign FP_adder_13ccs_42_io_in_a = FP_multiplier_10ccs_42_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_42_io_in_b = FPReg_42_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_43_clock = clock;
  assign FP_adder_13ccs_43_reset = reset;
  assign FP_adder_13ccs_43_io_in_a = FP_multiplier_10ccs_43_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_43_io_in_b = FPReg_43_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_44_clock = clock;
  assign FP_adder_13ccs_44_reset = reset;
  assign FP_adder_13ccs_44_io_in_a = FP_multiplier_10ccs_44_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_44_io_in_b = FPReg_44_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_45_clock = clock;
  assign FP_adder_13ccs_45_reset = reset;
  assign FP_adder_13ccs_45_io_in_a = FP_multiplier_10ccs_45_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_45_io_in_b = FPReg_45_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_46_clock = clock;
  assign FP_adder_13ccs_46_reset = reset;
  assign FP_adder_13ccs_46_io_in_a = FP_multiplier_10ccs_46_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_46_io_in_b = FPReg_46_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_47_clock = clock;
  assign FP_adder_13ccs_47_reset = reset;
  assign FP_adder_13ccs_47_io_in_a = FP_multiplier_10ccs_47_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_47_io_in_b = FPReg_47_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_48_clock = clock;
  assign FP_adder_13ccs_48_reset = reset;
  assign FP_adder_13ccs_48_io_in_a = FP_multiplier_10ccs_48_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_48_io_in_b = FPReg_48_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_49_clock = clock;
  assign FP_adder_13ccs_49_reset = reset;
  assign FP_adder_13ccs_49_io_in_a = FP_multiplier_10ccs_49_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_49_io_in_b = FPReg_49_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_50_clock = clock;
  assign FP_adder_13ccs_50_reset = reset;
  assign FP_adder_13ccs_50_io_in_a = FP_multiplier_10ccs_50_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_50_io_in_b = FPReg_50_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_51_clock = clock;
  assign FP_adder_13ccs_51_reset = reset;
  assign FP_adder_13ccs_51_io_in_a = FP_multiplier_10ccs_51_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_51_io_in_b = FPReg_51_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_52_clock = clock;
  assign FP_adder_13ccs_52_reset = reset;
  assign FP_adder_13ccs_52_io_in_a = FP_multiplier_10ccs_52_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_52_io_in_b = FPReg_52_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_53_clock = clock;
  assign FP_adder_13ccs_53_reset = reset;
  assign FP_adder_13ccs_53_io_in_a = FP_multiplier_10ccs_53_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_53_io_in_b = FPReg_53_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_54_clock = clock;
  assign FP_adder_13ccs_54_reset = reset;
  assign FP_adder_13ccs_54_io_in_a = FP_multiplier_10ccs_54_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_54_io_in_b = FPReg_54_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_55_clock = clock;
  assign FP_adder_13ccs_55_reset = reset;
  assign FP_adder_13ccs_55_io_in_a = FP_multiplier_10ccs_55_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_55_io_in_b = FPReg_55_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_56_clock = clock;
  assign FP_adder_13ccs_56_reset = reset;
  assign FP_adder_13ccs_56_io_in_a = FP_multiplier_10ccs_56_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_56_io_in_b = FPReg_56_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_57_clock = clock;
  assign FP_adder_13ccs_57_reset = reset;
  assign FP_adder_13ccs_57_io_in_a = FP_multiplier_10ccs_57_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_57_io_in_b = FPReg_57_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_58_clock = clock;
  assign FP_adder_13ccs_58_reset = reset;
  assign FP_adder_13ccs_58_io_in_a = FP_multiplier_10ccs_58_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_58_io_in_b = FPReg_58_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_59_clock = clock;
  assign FP_adder_13ccs_59_reset = reset;
  assign FP_adder_13ccs_59_io_in_a = FP_multiplier_10ccs_59_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_59_io_in_b = FPReg_59_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_60_clock = clock;
  assign FP_adder_13ccs_60_reset = reset;
  assign FP_adder_13ccs_60_io_in_a = FP_multiplier_10ccs_60_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_60_io_in_b = FPReg_60_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_61_clock = clock;
  assign FP_adder_13ccs_61_reset = reset;
  assign FP_adder_13ccs_61_io_in_a = FP_multiplier_10ccs_61_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_61_io_in_b = FPReg_61_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_62_clock = clock;
  assign FP_adder_13ccs_62_reset = reset;
  assign FP_adder_13ccs_62_io_in_a = FP_multiplier_10ccs_62_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_62_io_in_b = FPReg_62_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FP_adder_13ccs_63_clock = clock;
  assign FP_adder_13ccs_63_reset = reset;
  assign FP_adder_13ccs_63_io_in_a = FP_multiplier_10ccs_63_io_out_s; // @[FloatingPointDesigns.scala 2499:27]
  assign FP_adder_13ccs_63_io_in_b = FPReg_63_io_out; // @[FloatingPointDesigns.scala 2500:27]
  assign FPReg_clock = clock;
  assign FPReg_reset = reset;
  assign FPReg_io_in = io_in_c_0; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_1_clock = clock;
  assign FPReg_1_reset = reset;
  assign FPReg_1_io_in = io_in_c_1; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_2_clock = clock;
  assign FPReg_2_reset = reset;
  assign FPReg_2_io_in = io_in_c_2; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_3_clock = clock;
  assign FPReg_3_reset = reset;
  assign FPReg_3_io_in = io_in_c_3; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_4_clock = clock;
  assign FPReg_4_reset = reset;
  assign FPReg_4_io_in = io_in_c_4; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_5_clock = clock;
  assign FPReg_5_reset = reset;
  assign FPReg_5_io_in = io_in_c_5; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_6_clock = clock;
  assign FPReg_6_reset = reset;
  assign FPReg_6_io_in = io_in_c_6; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_7_clock = clock;
  assign FPReg_7_reset = reset;
  assign FPReg_7_io_in = io_in_c_7; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_8_clock = clock;
  assign FPReg_8_reset = reset;
  assign FPReg_8_io_in = io_in_c_8; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_9_clock = clock;
  assign FPReg_9_reset = reset;
  assign FPReg_9_io_in = io_in_c_9; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_10_clock = clock;
  assign FPReg_10_reset = reset;
  assign FPReg_10_io_in = io_in_c_10; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_11_clock = clock;
  assign FPReg_11_reset = reset;
  assign FPReg_11_io_in = io_in_c_11; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_12_clock = clock;
  assign FPReg_12_reset = reset;
  assign FPReg_12_io_in = io_in_c_12; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_13_clock = clock;
  assign FPReg_13_reset = reset;
  assign FPReg_13_io_in = io_in_c_13; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_14_clock = clock;
  assign FPReg_14_reset = reset;
  assign FPReg_14_io_in = io_in_c_14; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_15_clock = clock;
  assign FPReg_15_reset = reset;
  assign FPReg_15_io_in = io_in_c_15; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_16_clock = clock;
  assign FPReg_16_reset = reset;
  assign FPReg_16_io_in = io_in_c_16; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_17_clock = clock;
  assign FPReg_17_reset = reset;
  assign FPReg_17_io_in = io_in_c_17; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_18_clock = clock;
  assign FPReg_18_reset = reset;
  assign FPReg_18_io_in = io_in_c_18; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_19_clock = clock;
  assign FPReg_19_reset = reset;
  assign FPReg_19_io_in = io_in_c_19; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_20_clock = clock;
  assign FPReg_20_reset = reset;
  assign FPReg_20_io_in = io_in_c_20; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_21_clock = clock;
  assign FPReg_21_reset = reset;
  assign FPReg_21_io_in = io_in_c_21; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_22_clock = clock;
  assign FPReg_22_reset = reset;
  assign FPReg_22_io_in = io_in_c_22; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_23_clock = clock;
  assign FPReg_23_reset = reset;
  assign FPReg_23_io_in = io_in_c_23; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_24_clock = clock;
  assign FPReg_24_reset = reset;
  assign FPReg_24_io_in = io_in_c_24; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_25_clock = clock;
  assign FPReg_25_reset = reset;
  assign FPReg_25_io_in = io_in_c_25; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_26_clock = clock;
  assign FPReg_26_reset = reset;
  assign FPReg_26_io_in = io_in_c_26; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_27_clock = clock;
  assign FPReg_27_reset = reset;
  assign FPReg_27_io_in = io_in_c_27; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_28_clock = clock;
  assign FPReg_28_reset = reset;
  assign FPReg_28_io_in = io_in_c_28; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_29_clock = clock;
  assign FPReg_29_reset = reset;
  assign FPReg_29_io_in = io_in_c_29; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_30_clock = clock;
  assign FPReg_30_reset = reset;
  assign FPReg_30_io_in = io_in_c_30; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_31_clock = clock;
  assign FPReg_31_reset = reset;
  assign FPReg_31_io_in = io_in_c_31; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_32_clock = clock;
  assign FPReg_32_reset = reset;
  assign FPReg_32_io_in = io_in_c_32; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_33_clock = clock;
  assign FPReg_33_reset = reset;
  assign FPReg_33_io_in = io_in_c_33; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_34_clock = clock;
  assign FPReg_34_reset = reset;
  assign FPReg_34_io_in = io_in_c_34; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_35_clock = clock;
  assign FPReg_35_reset = reset;
  assign FPReg_35_io_in = io_in_c_35; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_36_clock = clock;
  assign FPReg_36_reset = reset;
  assign FPReg_36_io_in = io_in_c_36; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_37_clock = clock;
  assign FPReg_37_reset = reset;
  assign FPReg_37_io_in = io_in_c_37; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_38_clock = clock;
  assign FPReg_38_reset = reset;
  assign FPReg_38_io_in = io_in_c_38; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_39_clock = clock;
  assign FPReg_39_reset = reset;
  assign FPReg_39_io_in = io_in_c_39; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_40_clock = clock;
  assign FPReg_40_reset = reset;
  assign FPReg_40_io_in = io_in_c_40; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_41_clock = clock;
  assign FPReg_41_reset = reset;
  assign FPReg_41_io_in = io_in_c_41; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_42_clock = clock;
  assign FPReg_42_reset = reset;
  assign FPReg_42_io_in = io_in_c_42; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_43_clock = clock;
  assign FPReg_43_reset = reset;
  assign FPReg_43_io_in = io_in_c_43; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_44_clock = clock;
  assign FPReg_44_reset = reset;
  assign FPReg_44_io_in = io_in_c_44; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_45_clock = clock;
  assign FPReg_45_reset = reset;
  assign FPReg_45_io_in = io_in_c_45; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_46_clock = clock;
  assign FPReg_46_reset = reset;
  assign FPReg_46_io_in = io_in_c_46; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_47_clock = clock;
  assign FPReg_47_reset = reset;
  assign FPReg_47_io_in = io_in_c_47; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_48_clock = clock;
  assign FPReg_48_reset = reset;
  assign FPReg_48_io_in = io_in_c_48; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_49_clock = clock;
  assign FPReg_49_reset = reset;
  assign FPReg_49_io_in = io_in_c_49; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_50_clock = clock;
  assign FPReg_50_reset = reset;
  assign FPReg_50_io_in = io_in_c_50; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_51_clock = clock;
  assign FPReg_51_reset = reset;
  assign FPReg_51_io_in = io_in_c_51; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_52_clock = clock;
  assign FPReg_52_reset = reset;
  assign FPReg_52_io_in = io_in_c_52; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_53_clock = clock;
  assign FPReg_53_reset = reset;
  assign FPReg_53_io_in = io_in_c_53; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_54_clock = clock;
  assign FPReg_54_reset = reset;
  assign FPReg_54_io_in = io_in_c_54; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_55_clock = clock;
  assign FPReg_55_reset = reset;
  assign FPReg_55_io_in = io_in_c_55; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_56_clock = clock;
  assign FPReg_56_reset = reset;
  assign FPReg_56_io_in = io_in_c_56; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_57_clock = clock;
  assign FPReg_57_reset = reset;
  assign FPReg_57_io_in = io_in_c_57; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_58_clock = clock;
  assign FPReg_58_reset = reset;
  assign FPReg_58_io_in = io_in_c_58; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_59_clock = clock;
  assign FPReg_59_reset = reset;
  assign FPReg_59_io_in = io_in_c_59; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_60_clock = clock;
  assign FPReg_60_reset = reset;
  assign FPReg_60_io_in = io_in_c_60; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_61_clock = clock;
  assign FPReg_61_reset = reset;
  assign FPReg_61_io_in = io_in_c_61; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_62_clock = clock;
  assign FPReg_62_reset = reset;
  assign FPReg_62_io_in = io_in_c_62; // @[FloatingPointDesigns.scala 2498:25]
  assign FPReg_63_clock = clock;
  assign FPReg_63_reset = reset;
  assign FPReg_63_io_in = io_in_c_63; // @[FloatingPointDesigns.scala 2498:25]
endmodule
module hh_datapath_1(
  input           io_clk,
  input           io_rst,
  input  [15:0]   io_hh_cnt,
  input           io_d1_rdy,
  input           io_d1_vld,
  input           io_d2_vld,
  input           io_vk1_vld,
  input           io_d3_rdy,
  input           io_d3_vld,
  input           io_tk_vld,
  input           io_d4_rdy,
  input           io_d5_rdy,
  input           io_d5_vld,
  input           io_yj_sft,
  input           io_d4_sft,
  input  [2047:0] io_hh_din,
  output [2047:0] io_hh_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [2047:0] _RAND_0;
  reg [116223:0] _RAND_1;
  reg [116223:0] _RAND_2;
  reg [116223:0] _RAND_3;
  reg [116223:0] _RAND_4;
  reg [2047:0] _RAND_5;
  reg [2047:0] _RAND_6;
  reg [2047:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [4063:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
`endif // RANDOMIZE_REG_INIT
  wire  FP_DDOT_dp_clock; // @[hh_datapath_chisel.scala 248:21]
  wire  FP_DDOT_dp_reset; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_0; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_1; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_2; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_3; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_4; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_5; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_6; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_7; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_8; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_9; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_10; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_11; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_12; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_13; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_14; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_15; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_16; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_17; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_18; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_19; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_20; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_21; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_22; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_23; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_24; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_25; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_26; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_27; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_28; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_29; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_30; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_31; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_32; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_33; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_34; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_35; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_36; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_37; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_38; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_39; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_40; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_41; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_42; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_43; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_44; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_45; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_46; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_47; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_48; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_49; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_50; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_51; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_52; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_53; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_54; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_55; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_56; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_57; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_58; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_59; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_60; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_61; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_62; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_a_63; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_0; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_1; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_2; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_3; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_4; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_5; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_6; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_7; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_8; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_9; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_10; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_11; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_12; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_13; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_14; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_15; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_16; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_17; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_18; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_19; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_20; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_21; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_22; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_23; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_24; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_25; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_26; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_27; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_28; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_29; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_30; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_31; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_32; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_33; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_34; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_35; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_36; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_37; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_38; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_39; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_40; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_41; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_42; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_43; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_44; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_45; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_46; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_47; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_48; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_49; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_50; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_51; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_52; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_53; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_54; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_55; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_56; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_57; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_58; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_59; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_60; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_61; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_62; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_in_b_63; // @[hh_datapath_chisel.scala 248:21]
  wire [31:0] FP_DDOT_dp_io_out_s; // @[hh_datapath_chisel.scala 248:21]
  wire  FP_square_root_newfpu_clock; // @[hh_datapath_chisel.scala 256:22]
  wire  FP_square_root_newfpu_reset; // @[hh_datapath_chisel.scala 256:22]
  wire [31:0] FP_square_root_newfpu_io_in_a; // @[hh_datapath_chisel.scala 256:22]
  wire [31:0] FP_square_root_newfpu_io_out_s; // @[hh_datapath_chisel.scala 256:22]
  wire  hqr5_clock; // @[hh_datapath_chisel.scala 261:20]
  wire  hqr5_reset; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_in_a; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_in_b; // @[hh_datapath_chisel.scala 261:20]
  wire [31:0] hqr5_io_out_s; // @[hh_datapath_chisel.scala 261:20]
  wire  hqr7_clock; // @[hh_datapath_chisel.scala 266:20]
  wire  hqr7_reset; // @[hh_datapath_chisel.scala 266:20]
  wire [31:0] hqr7_io_in_a; // @[hh_datapath_chisel.scala 266:20]
  wire [31:0] hqr7_io_out_s; // @[hh_datapath_chisel.scala 266:20]
  wire  FP_multiplier_10ccs_clock; // @[hh_datapath_chisel.scala 270:21]
  wire  FP_multiplier_10ccs_reset; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_in_a; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_in_b; // @[hh_datapath_chisel.scala 270:21]
  wire [31:0] FP_multiplier_10ccs_io_out_s; // @[hh_datapath_chisel.scala 270:21]
  wire  axpy_dp_clock; // @[hh_datapath_chisel.scala 276:20]
  wire  axpy_dp_reset; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_a; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_b_63; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_in_c_63; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_0; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_1; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_2; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_3; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_4; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_5; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_6; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_7; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_8; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_9; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_10; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_11; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_12; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_13; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_14; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_15; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_16; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_17; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_18; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_19; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_20; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_21; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_22; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_23; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_24; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_25; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_26; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_27; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_28; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_29; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_30; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_31; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_32; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_33; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_34; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_35; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_36; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_37; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_38; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_39; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_40; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_41; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_42; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_43; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_44; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_45; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_46; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_47; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_48; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_49; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_50; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_51; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_52; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_53; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_54; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_55; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_56; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_57; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_58; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_59; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_60; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_61; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_62; // @[hh_datapath_chisel.scala 276:20]
  wire [31:0] axpy_dp_io_out_s_63; // @[hh_datapath_chisel.scala 276:20]
  reg [2047:0] yj0; // @[hh_datapath_chisel.scala 53:18]
  reg [116223:0] yj_reg_1; // @[hh_datapath_chisel.scala 54:23]
  reg [116223:0] yj_reg_2; // @[hh_datapath_chisel.scala 55:23]
  reg [116223:0] yj_reg_3; // @[hh_datapath_chisel.scala 56:23]
  reg [116223:0] yj_reg_4; // @[hh_datapath_chisel.scala 57:23]
  wire [118271:0] _yj_reg_4_T_1 = {yj_reg_3[2047:0],yj_reg_4}; // @[Cat.scala 31:58]
  wire [118271:0] _yj_reg_3_T_1 = {yj_reg_2[2047:0],yj_reg_3}; // @[Cat.scala 31:58]
  wire [118271:0] _yj_reg_2_T_1 = {yj_reg_1[2047:0],yj_reg_2}; // @[Cat.scala 31:58]
  wire [118271:0] _yj_reg_1_T = {io_hh_din,yj_reg_1}; // @[Cat.scala 31:58]
  reg [2047:0] ddot_din_a_reg; // @[hh_datapath_chisel.scala 82:29]
  reg [2047:0] ddot_din_b_reg; // @[hh_datapath_chisel.scala 83:29]
  reg [2047:0] vk_reg; // @[hh_datapath_chisel.scala 85:21]
  reg [31:0] d1_reg; // @[hh_datapath_chisel.scala 86:21]
  reg [31:0] d3_reg; // @[hh_datapath_chisel.scala 87:21]
  reg [31:0] d4_update; // @[hh_datapath_chisel.scala 93:24]
  reg [31:0] x1_reg; // @[hh_datapath_chisel.scala 102:21]
  reg [31:0] d2_reg; // @[hh_datapath_chisel.scala 103:21]
  reg [31:0] vk1_reg; // @[hh_datapath_chisel.scala 104:22]
  reg [31:0] tk_reg; // @[hh_datapath_chisel.scala 105:21]
  reg [31:0] d4_reg; // @[hh_datapath_chisel.scala 106:21]
  reg [31:0] d5_reg; // @[hh_datapath_chisel.scala 107:21]
  wire [31:0] vk1_update = hqr5_io_out_s; // @[hh_datapath_chisel.scala 264:15 91:26]
  wire [31:0] vk1 = io_vk1_vld ? vk1_update : vk1_reg; // @[hh_datapath_chisel.scala 195:21 196:11 198:11]
  wire [15:0] _myNewVec_63_T_1 = io_hh_cnt + 16'h1; // @[hh_datapath_chisel.scala 234:55]
  wire [16:0] _myNewVec_63_T_2 = {{1'd0}, _myNewVec_63_T_1}; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] myVec_63 = io_hh_din[31:0]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_62 = io_hh_din[63:32]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_61 = io_hh_din[95:64]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_60 = io_hh_din[127:96]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_59 = io_hh_din[159:128]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_58 = io_hh_din[191:160]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_57 = io_hh_din[223:192]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_56 = io_hh_din[255:224]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_55 = io_hh_din[287:256]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_54 = io_hh_din[319:288]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_53 = io_hh_din[351:320]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_52 = io_hh_din[383:352]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_51 = io_hh_din[415:384]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_50 = io_hh_din[447:416]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_49 = io_hh_din[479:448]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_48 = io_hh_din[511:480]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_47 = io_hh_din[543:512]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_46 = io_hh_din[575:544]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_45 = io_hh_din[607:576]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_44 = io_hh_din[639:608]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_43 = io_hh_din[671:640]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_42 = io_hh_din[703:672]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_41 = io_hh_din[735:704]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_40 = io_hh_din[767:736]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_39 = io_hh_din[799:768]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_38 = io_hh_din[831:800]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_37 = io_hh_din[863:832]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_36 = io_hh_din[895:864]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_35 = io_hh_din[927:896]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_34 = io_hh_din[959:928]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_33 = io_hh_din[991:960]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_32 = io_hh_din[1023:992]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_31 = io_hh_din[1055:1024]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_30 = io_hh_din[1087:1056]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_29 = io_hh_din[1119:1088]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_28 = io_hh_din[1151:1120]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_27 = io_hh_din[1183:1152]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_26 = io_hh_din[1215:1184]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_25 = io_hh_din[1247:1216]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_24 = io_hh_din[1279:1248]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_23 = io_hh_din[1311:1280]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_22 = io_hh_din[1343:1312]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_21 = io_hh_din[1375:1344]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_20 = io_hh_din[1407:1376]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_19 = io_hh_din[1439:1408]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_18 = io_hh_din[1471:1440]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_17 = io_hh_din[1503:1472]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_16 = io_hh_din[1535:1504]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_15 = io_hh_din[1567:1536]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_14 = io_hh_din[1599:1568]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_13 = io_hh_din[1631:1600]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_12 = io_hh_din[1663:1632]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_11 = io_hh_din[1695:1664]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_10 = io_hh_din[1727:1696]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_9 = io_hh_din[1759:1728]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_8 = io_hh_din[1791:1760]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_7 = io_hh_din[1823:1792]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_6 = io_hh_din[1855:1824]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_5 = io_hh_din[1887:1856]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_4 = io_hh_din[1919:1888]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_3 = io_hh_din[1951:1920]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_2 = io_hh_din[1983:1952]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_1 = io_hh_din[2015:1984]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] myVec_0 = io_hh_din[2047:2016]; // @[hh_datapath_chisel.scala 221:28]
  wire [31:0] _GEN_107 = 6'h1 == _myNewVec_63_T_2[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_108 = 6'h2 == _myNewVec_63_T_2[5:0] ? myVec_2 : _GEN_107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_109 = 6'h3 == _myNewVec_63_T_2[5:0] ? myVec_3 : _GEN_108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_110 = 6'h4 == _myNewVec_63_T_2[5:0] ? myVec_4 : _GEN_109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_111 = 6'h5 == _myNewVec_63_T_2[5:0] ? myVec_5 : _GEN_110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_112 = 6'h6 == _myNewVec_63_T_2[5:0] ? myVec_6 : _GEN_111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_113 = 6'h7 == _myNewVec_63_T_2[5:0] ? myVec_7 : _GEN_112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_114 = 6'h8 == _myNewVec_63_T_2[5:0] ? myVec_8 : _GEN_113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_115 = 6'h9 == _myNewVec_63_T_2[5:0] ? myVec_9 : _GEN_114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_116 = 6'ha == _myNewVec_63_T_2[5:0] ? myVec_10 : _GEN_115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_117 = 6'hb == _myNewVec_63_T_2[5:0] ? myVec_11 : _GEN_116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_118 = 6'hc == _myNewVec_63_T_2[5:0] ? myVec_12 : _GEN_117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_119 = 6'hd == _myNewVec_63_T_2[5:0] ? myVec_13 : _GEN_118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_120 = 6'he == _myNewVec_63_T_2[5:0] ? myVec_14 : _GEN_119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_121 = 6'hf == _myNewVec_63_T_2[5:0] ? myVec_15 : _GEN_120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_122 = 6'h10 == _myNewVec_63_T_2[5:0] ? myVec_16 : _GEN_121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_123 = 6'h11 == _myNewVec_63_T_2[5:0] ? myVec_17 : _GEN_122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_124 = 6'h12 == _myNewVec_63_T_2[5:0] ? myVec_18 : _GEN_123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_125 = 6'h13 == _myNewVec_63_T_2[5:0] ? myVec_19 : _GEN_124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_126 = 6'h14 == _myNewVec_63_T_2[5:0] ? myVec_20 : _GEN_125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_127 = 6'h15 == _myNewVec_63_T_2[5:0] ? myVec_21 : _GEN_126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_128 = 6'h16 == _myNewVec_63_T_2[5:0] ? myVec_22 : _GEN_127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_129 = 6'h17 == _myNewVec_63_T_2[5:0] ? myVec_23 : _GEN_128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_130 = 6'h18 == _myNewVec_63_T_2[5:0] ? myVec_24 : _GEN_129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_131 = 6'h19 == _myNewVec_63_T_2[5:0] ? myVec_25 : _GEN_130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_132 = 6'h1a == _myNewVec_63_T_2[5:0] ? myVec_26 : _GEN_131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_133 = 6'h1b == _myNewVec_63_T_2[5:0] ? myVec_27 : _GEN_132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_134 = 6'h1c == _myNewVec_63_T_2[5:0] ? myVec_28 : _GEN_133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_135 = 6'h1d == _myNewVec_63_T_2[5:0] ? myVec_29 : _GEN_134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_136 = 6'h1e == _myNewVec_63_T_2[5:0] ? myVec_30 : _GEN_135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_137 = 6'h1f == _myNewVec_63_T_2[5:0] ? myVec_31 : _GEN_136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_138 = 6'h20 == _myNewVec_63_T_2[5:0] ? myVec_32 : _GEN_137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_139 = 6'h21 == _myNewVec_63_T_2[5:0] ? myVec_33 : _GEN_138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_140 = 6'h22 == _myNewVec_63_T_2[5:0] ? myVec_34 : _GEN_139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_141 = 6'h23 == _myNewVec_63_T_2[5:0] ? myVec_35 : _GEN_140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_142 = 6'h24 == _myNewVec_63_T_2[5:0] ? myVec_36 : _GEN_141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_143 = 6'h25 == _myNewVec_63_T_2[5:0] ? myVec_37 : _GEN_142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_144 = 6'h26 == _myNewVec_63_T_2[5:0] ? myVec_38 : _GEN_143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_145 = 6'h27 == _myNewVec_63_T_2[5:0] ? myVec_39 : _GEN_144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_146 = 6'h28 == _myNewVec_63_T_2[5:0] ? myVec_40 : _GEN_145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_147 = 6'h29 == _myNewVec_63_T_2[5:0] ? myVec_41 : _GEN_146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_148 = 6'h2a == _myNewVec_63_T_2[5:0] ? myVec_42 : _GEN_147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_149 = 6'h2b == _myNewVec_63_T_2[5:0] ? myVec_43 : _GEN_148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_150 = 6'h2c == _myNewVec_63_T_2[5:0] ? myVec_44 : _GEN_149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_151 = 6'h2d == _myNewVec_63_T_2[5:0] ? myVec_45 : _GEN_150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_152 = 6'h2e == _myNewVec_63_T_2[5:0] ? myVec_46 : _GEN_151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_153 = 6'h2f == _myNewVec_63_T_2[5:0] ? myVec_47 : _GEN_152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_154 = 6'h30 == _myNewVec_63_T_2[5:0] ? myVec_48 : _GEN_153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_155 = 6'h31 == _myNewVec_63_T_2[5:0] ? myVec_49 : _GEN_154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_156 = 6'h32 == _myNewVec_63_T_2[5:0] ? myVec_50 : _GEN_155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_157 = 6'h33 == _myNewVec_63_T_2[5:0] ? myVec_51 : _GEN_156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_158 = 6'h34 == _myNewVec_63_T_2[5:0] ? myVec_52 : _GEN_157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_159 = 6'h35 == _myNewVec_63_T_2[5:0] ? myVec_53 : _GEN_158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_160 = 6'h36 == _myNewVec_63_T_2[5:0] ? myVec_54 : _GEN_159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_161 = 6'h37 == _myNewVec_63_T_2[5:0] ? myVec_55 : _GEN_160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_162 = 6'h38 == _myNewVec_63_T_2[5:0] ? myVec_56 : _GEN_161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_163 = 6'h39 == _myNewVec_63_T_2[5:0] ? myVec_57 : _GEN_162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_164 = 6'h3a == _myNewVec_63_T_2[5:0] ? myVec_58 : _GEN_163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_165 = 6'h3b == _myNewVec_63_T_2[5:0] ? myVec_59 : _GEN_164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_166 = 6'h3c == _myNewVec_63_T_2[5:0] ? myVec_60 : _GEN_165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_167 = 6'h3d == _myNewVec_63_T_2[5:0] ? myVec_61 : _GEN_166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_168 = 6'h3e == _myNewVec_63_T_2[5:0] ? myVec_62 : _GEN_167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_63 = 6'h3f == _myNewVec_63_T_2[5:0] ? myVec_63 : _GEN_168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_62_T_3 = _myNewVec_63_T_1 + 16'h1; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_171 = 6'h1 == _myNewVec_62_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_172 = 6'h2 == _myNewVec_62_T_3[5:0] ? myVec_2 : _GEN_171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_173 = 6'h3 == _myNewVec_62_T_3[5:0] ? myVec_3 : _GEN_172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_174 = 6'h4 == _myNewVec_62_T_3[5:0] ? myVec_4 : _GEN_173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_175 = 6'h5 == _myNewVec_62_T_3[5:0] ? myVec_5 : _GEN_174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_176 = 6'h6 == _myNewVec_62_T_3[5:0] ? myVec_6 : _GEN_175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_177 = 6'h7 == _myNewVec_62_T_3[5:0] ? myVec_7 : _GEN_176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_178 = 6'h8 == _myNewVec_62_T_3[5:0] ? myVec_8 : _GEN_177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_179 = 6'h9 == _myNewVec_62_T_3[5:0] ? myVec_9 : _GEN_178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_180 = 6'ha == _myNewVec_62_T_3[5:0] ? myVec_10 : _GEN_179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_181 = 6'hb == _myNewVec_62_T_3[5:0] ? myVec_11 : _GEN_180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_182 = 6'hc == _myNewVec_62_T_3[5:0] ? myVec_12 : _GEN_181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_183 = 6'hd == _myNewVec_62_T_3[5:0] ? myVec_13 : _GEN_182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_184 = 6'he == _myNewVec_62_T_3[5:0] ? myVec_14 : _GEN_183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_185 = 6'hf == _myNewVec_62_T_3[5:0] ? myVec_15 : _GEN_184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_186 = 6'h10 == _myNewVec_62_T_3[5:0] ? myVec_16 : _GEN_185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_187 = 6'h11 == _myNewVec_62_T_3[5:0] ? myVec_17 : _GEN_186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_188 = 6'h12 == _myNewVec_62_T_3[5:0] ? myVec_18 : _GEN_187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_189 = 6'h13 == _myNewVec_62_T_3[5:0] ? myVec_19 : _GEN_188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_190 = 6'h14 == _myNewVec_62_T_3[5:0] ? myVec_20 : _GEN_189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_191 = 6'h15 == _myNewVec_62_T_3[5:0] ? myVec_21 : _GEN_190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_192 = 6'h16 == _myNewVec_62_T_3[5:0] ? myVec_22 : _GEN_191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_193 = 6'h17 == _myNewVec_62_T_3[5:0] ? myVec_23 : _GEN_192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_194 = 6'h18 == _myNewVec_62_T_3[5:0] ? myVec_24 : _GEN_193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_195 = 6'h19 == _myNewVec_62_T_3[5:0] ? myVec_25 : _GEN_194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_196 = 6'h1a == _myNewVec_62_T_3[5:0] ? myVec_26 : _GEN_195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_197 = 6'h1b == _myNewVec_62_T_3[5:0] ? myVec_27 : _GEN_196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_198 = 6'h1c == _myNewVec_62_T_3[5:0] ? myVec_28 : _GEN_197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_199 = 6'h1d == _myNewVec_62_T_3[5:0] ? myVec_29 : _GEN_198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_200 = 6'h1e == _myNewVec_62_T_3[5:0] ? myVec_30 : _GEN_199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_201 = 6'h1f == _myNewVec_62_T_3[5:0] ? myVec_31 : _GEN_200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_202 = 6'h20 == _myNewVec_62_T_3[5:0] ? myVec_32 : _GEN_201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_203 = 6'h21 == _myNewVec_62_T_3[5:0] ? myVec_33 : _GEN_202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_204 = 6'h22 == _myNewVec_62_T_3[5:0] ? myVec_34 : _GEN_203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_205 = 6'h23 == _myNewVec_62_T_3[5:0] ? myVec_35 : _GEN_204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_206 = 6'h24 == _myNewVec_62_T_3[5:0] ? myVec_36 : _GEN_205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_207 = 6'h25 == _myNewVec_62_T_3[5:0] ? myVec_37 : _GEN_206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_208 = 6'h26 == _myNewVec_62_T_3[5:0] ? myVec_38 : _GEN_207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_209 = 6'h27 == _myNewVec_62_T_3[5:0] ? myVec_39 : _GEN_208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_210 = 6'h28 == _myNewVec_62_T_3[5:0] ? myVec_40 : _GEN_209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_211 = 6'h29 == _myNewVec_62_T_3[5:0] ? myVec_41 : _GEN_210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_212 = 6'h2a == _myNewVec_62_T_3[5:0] ? myVec_42 : _GEN_211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_213 = 6'h2b == _myNewVec_62_T_3[5:0] ? myVec_43 : _GEN_212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_214 = 6'h2c == _myNewVec_62_T_3[5:0] ? myVec_44 : _GEN_213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_215 = 6'h2d == _myNewVec_62_T_3[5:0] ? myVec_45 : _GEN_214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_216 = 6'h2e == _myNewVec_62_T_3[5:0] ? myVec_46 : _GEN_215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_217 = 6'h2f == _myNewVec_62_T_3[5:0] ? myVec_47 : _GEN_216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_218 = 6'h30 == _myNewVec_62_T_3[5:0] ? myVec_48 : _GEN_217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_219 = 6'h31 == _myNewVec_62_T_3[5:0] ? myVec_49 : _GEN_218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_220 = 6'h32 == _myNewVec_62_T_3[5:0] ? myVec_50 : _GEN_219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_221 = 6'h33 == _myNewVec_62_T_3[5:0] ? myVec_51 : _GEN_220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_222 = 6'h34 == _myNewVec_62_T_3[5:0] ? myVec_52 : _GEN_221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_223 = 6'h35 == _myNewVec_62_T_3[5:0] ? myVec_53 : _GEN_222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_224 = 6'h36 == _myNewVec_62_T_3[5:0] ? myVec_54 : _GEN_223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_225 = 6'h37 == _myNewVec_62_T_3[5:0] ? myVec_55 : _GEN_224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_226 = 6'h38 == _myNewVec_62_T_3[5:0] ? myVec_56 : _GEN_225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_227 = 6'h39 == _myNewVec_62_T_3[5:0] ? myVec_57 : _GEN_226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_228 = 6'h3a == _myNewVec_62_T_3[5:0] ? myVec_58 : _GEN_227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_229 = 6'h3b == _myNewVec_62_T_3[5:0] ? myVec_59 : _GEN_228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_230 = 6'h3c == _myNewVec_62_T_3[5:0] ? myVec_60 : _GEN_229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_231 = 6'h3d == _myNewVec_62_T_3[5:0] ? myVec_61 : _GEN_230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_232 = 6'h3e == _myNewVec_62_T_3[5:0] ? myVec_62 : _GEN_231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_62 = 6'h3f == _myNewVec_62_T_3[5:0] ? myVec_63 : _GEN_232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_61_T_3 = _myNewVec_63_T_1 + 16'h2; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_235 = 6'h1 == _myNewVec_61_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_236 = 6'h2 == _myNewVec_61_T_3[5:0] ? myVec_2 : _GEN_235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_237 = 6'h3 == _myNewVec_61_T_3[5:0] ? myVec_3 : _GEN_236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_238 = 6'h4 == _myNewVec_61_T_3[5:0] ? myVec_4 : _GEN_237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_239 = 6'h5 == _myNewVec_61_T_3[5:0] ? myVec_5 : _GEN_238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_240 = 6'h6 == _myNewVec_61_T_3[5:0] ? myVec_6 : _GEN_239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_241 = 6'h7 == _myNewVec_61_T_3[5:0] ? myVec_7 : _GEN_240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_242 = 6'h8 == _myNewVec_61_T_3[5:0] ? myVec_8 : _GEN_241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_243 = 6'h9 == _myNewVec_61_T_3[5:0] ? myVec_9 : _GEN_242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_244 = 6'ha == _myNewVec_61_T_3[5:0] ? myVec_10 : _GEN_243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_245 = 6'hb == _myNewVec_61_T_3[5:0] ? myVec_11 : _GEN_244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_246 = 6'hc == _myNewVec_61_T_3[5:0] ? myVec_12 : _GEN_245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_247 = 6'hd == _myNewVec_61_T_3[5:0] ? myVec_13 : _GEN_246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_248 = 6'he == _myNewVec_61_T_3[5:0] ? myVec_14 : _GEN_247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_249 = 6'hf == _myNewVec_61_T_3[5:0] ? myVec_15 : _GEN_248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_250 = 6'h10 == _myNewVec_61_T_3[5:0] ? myVec_16 : _GEN_249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_251 = 6'h11 == _myNewVec_61_T_3[5:0] ? myVec_17 : _GEN_250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_252 = 6'h12 == _myNewVec_61_T_3[5:0] ? myVec_18 : _GEN_251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_253 = 6'h13 == _myNewVec_61_T_3[5:0] ? myVec_19 : _GEN_252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_254 = 6'h14 == _myNewVec_61_T_3[5:0] ? myVec_20 : _GEN_253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_255 = 6'h15 == _myNewVec_61_T_3[5:0] ? myVec_21 : _GEN_254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_256 = 6'h16 == _myNewVec_61_T_3[5:0] ? myVec_22 : _GEN_255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_257 = 6'h17 == _myNewVec_61_T_3[5:0] ? myVec_23 : _GEN_256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_258 = 6'h18 == _myNewVec_61_T_3[5:0] ? myVec_24 : _GEN_257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_259 = 6'h19 == _myNewVec_61_T_3[5:0] ? myVec_25 : _GEN_258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_260 = 6'h1a == _myNewVec_61_T_3[5:0] ? myVec_26 : _GEN_259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_261 = 6'h1b == _myNewVec_61_T_3[5:0] ? myVec_27 : _GEN_260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_262 = 6'h1c == _myNewVec_61_T_3[5:0] ? myVec_28 : _GEN_261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_263 = 6'h1d == _myNewVec_61_T_3[5:0] ? myVec_29 : _GEN_262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_264 = 6'h1e == _myNewVec_61_T_3[5:0] ? myVec_30 : _GEN_263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_265 = 6'h1f == _myNewVec_61_T_3[5:0] ? myVec_31 : _GEN_264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_266 = 6'h20 == _myNewVec_61_T_3[5:0] ? myVec_32 : _GEN_265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_267 = 6'h21 == _myNewVec_61_T_3[5:0] ? myVec_33 : _GEN_266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_268 = 6'h22 == _myNewVec_61_T_3[5:0] ? myVec_34 : _GEN_267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_269 = 6'h23 == _myNewVec_61_T_3[5:0] ? myVec_35 : _GEN_268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_270 = 6'h24 == _myNewVec_61_T_3[5:0] ? myVec_36 : _GEN_269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_271 = 6'h25 == _myNewVec_61_T_3[5:0] ? myVec_37 : _GEN_270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_272 = 6'h26 == _myNewVec_61_T_3[5:0] ? myVec_38 : _GEN_271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_273 = 6'h27 == _myNewVec_61_T_3[5:0] ? myVec_39 : _GEN_272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_274 = 6'h28 == _myNewVec_61_T_3[5:0] ? myVec_40 : _GEN_273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_275 = 6'h29 == _myNewVec_61_T_3[5:0] ? myVec_41 : _GEN_274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_276 = 6'h2a == _myNewVec_61_T_3[5:0] ? myVec_42 : _GEN_275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_277 = 6'h2b == _myNewVec_61_T_3[5:0] ? myVec_43 : _GEN_276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_278 = 6'h2c == _myNewVec_61_T_3[5:0] ? myVec_44 : _GEN_277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_279 = 6'h2d == _myNewVec_61_T_3[5:0] ? myVec_45 : _GEN_278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_280 = 6'h2e == _myNewVec_61_T_3[5:0] ? myVec_46 : _GEN_279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_281 = 6'h2f == _myNewVec_61_T_3[5:0] ? myVec_47 : _GEN_280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_282 = 6'h30 == _myNewVec_61_T_3[5:0] ? myVec_48 : _GEN_281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_283 = 6'h31 == _myNewVec_61_T_3[5:0] ? myVec_49 : _GEN_282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_284 = 6'h32 == _myNewVec_61_T_3[5:0] ? myVec_50 : _GEN_283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_285 = 6'h33 == _myNewVec_61_T_3[5:0] ? myVec_51 : _GEN_284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_286 = 6'h34 == _myNewVec_61_T_3[5:0] ? myVec_52 : _GEN_285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_287 = 6'h35 == _myNewVec_61_T_3[5:0] ? myVec_53 : _GEN_286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_288 = 6'h36 == _myNewVec_61_T_3[5:0] ? myVec_54 : _GEN_287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_289 = 6'h37 == _myNewVec_61_T_3[5:0] ? myVec_55 : _GEN_288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_290 = 6'h38 == _myNewVec_61_T_3[5:0] ? myVec_56 : _GEN_289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_291 = 6'h39 == _myNewVec_61_T_3[5:0] ? myVec_57 : _GEN_290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_292 = 6'h3a == _myNewVec_61_T_3[5:0] ? myVec_58 : _GEN_291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_293 = 6'h3b == _myNewVec_61_T_3[5:0] ? myVec_59 : _GEN_292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_294 = 6'h3c == _myNewVec_61_T_3[5:0] ? myVec_60 : _GEN_293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_295 = 6'h3d == _myNewVec_61_T_3[5:0] ? myVec_61 : _GEN_294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_296 = 6'h3e == _myNewVec_61_T_3[5:0] ? myVec_62 : _GEN_295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_61 = 6'h3f == _myNewVec_61_T_3[5:0] ? myVec_63 : _GEN_296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_60_T_3 = _myNewVec_63_T_1 + 16'h3; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_299 = 6'h1 == _myNewVec_60_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_300 = 6'h2 == _myNewVec_60_T_3[5:0] ? myVec_2 : _GEN_299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_301 = 6'h3 == _myNewVec_60_T_3[5:0] ? myVec_3 : _GEN_300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_302 = 6'h4 == _myNewVec_60_T_3[5:0] ? myVec_4 : _GEN_301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_303 = 6'h5 == _myNewVec_60_T_3[5:0] ? myVec_5 : _GEN_302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_304 = 6'h6 == _myNewVec_60_T_3[5:0] ? myVec_6 : _GEN_303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_305 = 6'h7 == _myNewVec_60_T_3[5:0] ? myVec_7 : _GEN_304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_306 = 6'h8 == _myNewVec_60_T_3[5:0] ? myVec_8 : _GEN_305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_307 = 6'h9 == _myNewVec_60_T_3[5:0] ? myVec_9 : _GEN_306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_308 = 6'ha == _myNewVec_60_T_3[5:0] ? myVec_10 : _GEN_307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_309 = 6'hb == _myNewVec_60_T_3[5:0] ? myVec_11 : _GEN_308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_310 = 6'hc == _myNewVec_60_T_3[5:0] ? myVec_12 : _GEN_309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_311 = 6'hd == _myNewVec_60_T_3[5:0] ? myVec_13 : _GEN_310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_312 = 6'he == _myNewVec_60_T_3[5:0] ? myVec_14 : _GEN_311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_313 = 6'hf == _myNewVec_60_T_3[5:0] ? myVec_15 : _GEN_312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_314 = 6'h10 == _myNewVec_60_T_3[5:0] ? myVec_16 : _GEN_313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_315 = 6'h11 == _myNewVec_60_T_3[5:0] ? myVec_17 : _GEN_314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_316 = 6'h12 == _myNewVec_60_T_3[5:0] ? myVec_18 : _GEN_315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_317 = 6'h13 == _myNewVec_60_T_3[5:0] ? myVec_19 : _GEN_316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_318 = 6'h14 == _myNewVec_60_T_3[5:0] ? myVec_20 : _GEN_317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_319 = 6'h15 == _myNewVec_60_T_3[5:0] ? myVec_21 : _GEN_318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_320 = 6'h16 == _myNewVec_60_T_3[5:0] ? myVec_22 : _GEN_319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_321 = 6'h17 == _myNewVec_60_T_3[5:0] ? myVec_23 : _GEN_320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_322 = 6'h18 == _myNewVec_60_T_3[5:0] ? myVec_24 : _GEN_321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_323 = 6'h19 == _myNewVec_60_T_3[5:0] ? myVec_25 : _GEN_322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_324 = 6'h1a == _myNewVec_60_T_3[5:0] ? myVec_26 : _GEN_323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_325 = 6'h1b == _myNewVec_60_T_3[5:0] ? myVec_27 : _GEN_324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_326 = 6'h1c == _myNewVec_60_T_3[5:0] ? myVec_28 : _GEN_325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_327 = 6'h1d == _myNewVec_60_T_3[5:0] ? myVec_29 : _GEN_326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_328 = 6'h1e == _myNewVec_60_T_3[5:0] ? myVec_30 : _GEN_327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_329 = 6'h1f == _myNewVec_60_T_3[5:0] ? myVec_31 : _GEN_328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_330 = 6'h20 == _myNewVec_60_T_3[5:0] ? myVec_32 : _GEN_329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_331 = 6'h21 == _myNewVec_60_T_3[5:0] ? myVec_33 : _GEN_330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_332 = 6'h22 == _myNewVec_60_T_3[5:0] ? myVec_34 : _GEN_331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_333 = 6'h23 == _myNewVec_60_T_3[5:0] ? myVec_35 : _GEN_332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_334 = 6'h24 == _myNewVec_60_T_3[5:0] ? myVec_36 : _GEN_333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_335 = 6'h25 == _myNewVec_60_T_3[5:0] ? myVec_37 : _GEN_334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_336 = 6'h26 == _myNewVec_60_T_3[5:0] ? myVec_38 : _GEN_335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_337 = 6'h27 == _myNewVec_60_T_3[5:0] ? myVec_39 : _GEN_336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_338 = 6'h28 == _myNewVec_60_T_3[5:0] ? myVec_40 : _GEN_337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_339 = 6'h29 == _myNewVec_60_T_3[5:0] ? myVec_41 : _GEN_338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_340 = 6'h2a == _myNewVec_60_T_3[5:0] ? myVec_42 : _GEN_339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_341 = 6'h2b == _myNewVec_60_T_3[5:0] ? myVec_43 : _GEN_340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_342 = 6'h2c == _myNewVec_60_T_3[5:0] ? myVec_44 : _GEN_341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_343 = 6'h2d == _myNewVec_60_T_3[5:0] ? myVec_45 : _GEN_342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_344 = 6'h2e == _myNewVec_60_T_3[5:0] ? myVec_46 : _GEN_343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_345 = 6'h2f == _myNewVec_60_T_3[5:0] ? myVec_47 : _GEN_344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_346 = 6'h30 == _myNewVec_60_T_3[5:0] ? myVec_48 : _GEN_345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_347 = 6'h31 == _myNewVec_60_T_3[5:0] ? myVec_49 : _GEN_346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_348 = 6'h32 == _myNewVec_60_T_3[5:0] ? myVec_50 : _GEN_347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_349 = 6'h33 == _myNewVec_60_T_3[5:0] ? myVec_51 : _GEN_348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_350 = 6'h34 == _myNewVec_60_T_3[5:0] ? myVec_52 : _GEN_349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_351 = 6'h35 == _myNewVec_60_T_3[5:0] ? myVec_53 : _GEN_350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_352 = 6'h36 == _myNewVec_60_T_3[5:0] ? myVec_54 : _GEN_351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_353 = 6'h37 == _myNewVec_60_T_3[5:0] ? myVec_55 : _GEN_352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_354 = 6'h38 == _myNewVec_60_T_3[5:0] ? myVec_56 : _GEN_353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_355 = 6'h39 == _myNewVec_60_T_3[5:0] ? myVec_57 : _GEN_354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_356 = 6'h3a == _myNewVec_60_T_3[5:0] ? myVec_58 : _GEN_355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_357 = 6'h3b == _myNewVec_60_T_3[5:0] ? myVec_59 : _GEN_356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_358 = 6'h3c == _myNewVec_60_T_3[5:0] ? myVec_60 : _GEN_357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_359 = 6'h3d == _myNewVec_60_T_3[5:0] ? myVec_61 : _GEN_358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_360 = 6'h3e == _myNewVec_60_T_3[5:0] ? myVec_62 : _GEN_359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_60 = 6'h3f == _myNewVec_60_T_3[5:0] ? myVec_63 : _GEN_360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_59_T_3 = _myNewVec_63_T_1 + 16'h4; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_363 = 6'h1 == _myNewVec_59_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_364 = 6'h2 == _myNewVec_59_T_3[5:0] ? myVec_2 : _GEN_363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_365 = 6'h3 == _myNewVec_59_T_3[5:0] ? myVec_3 : _GEN_364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_366 = 6'h4 == _myNewVec_59_T_3[5:0] ? myVec_4 : _GEN_365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_367 = 6'h5 == _myNewVec_59_T_3[5:0] ? myVec_5 : _GEN_366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_368 = 6'h6 == _myNewVec_59_T_3[5:0] ? myVec_6 : _GEN_367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_369 = 6'h7 == _myNewVec_59_T_3[5:0] ? myVec_7 : _GEN_368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_370 = 6'h8 == _myNewVec_59_T_3[5:0] ? myVec_8 : _GEN_369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_371 = 6'h9 == _myNewVec_59_T_3[5:0] ? myVec_9 : _GEN_370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_372 = 6'ha == _myNewVec_59_T_3[5:0] ? myVec_10 : _GEN_371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_373 = 6'hb == _myNewVec_59_T_3[5:0] ? myVec_11 : _GEN_372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_374 = 6'hc == _myNewVec_59_T_3[5:0] ? myVec_12 : _GEN_373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_375 = 6'hd == _myNewVec_59_T_3[5:0] ? myVec_13 : _GEN_374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_376 = 6'he == _myNewVec_59_T_3[5:0] ? myVec_14 : _GEN_375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_377 = 6'hf == _myNewVec_59_T_3[5:0] ? myVec_15 : _GEN_376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_378 = 6'h10 == _myNewVec_59_T_3[5:0] ? myVec_16 : _GEN_377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_379 = 6'h11 == _myNewVec_59_T_3[5:0] ? myVec_17 : _GEN_378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_380 = 6'h12 == _myNewVec_59_T_3[5:0] ? myVec_18 : _GEN_379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_381 = 6'h13 == _myNewVec_59_T_3[5:0] ? myVec_19 : _GEN_380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_382 = 6'h14 == _myNewVec_59_T_3[5:0] ? myVec_20 : _GEN_381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_383 = 6'h15 == _myNewVec_59_T_3[5:0] ? myVec_21 : _GEN_382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_384 = 6'h16 == _myNewVec_59_T_3[5:0] ? myVec_22 : _GEN_383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_385 = 6'h17 == _myNewVec_59_T_3[5:0] ? myVec_23 : _GEN_384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_386 = 6'h18 == _myNewVec_59_T_3[5:0] ? myVec_24 : _GEN_385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_387 = 6'h19 == _myNewVec_59_T_3[5:0] ? myVec_25 : _GEN_386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_388 = 6'h1a == _myNewVec_59_T_3[5:0] ? myVec_26 : _GEN_387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_389 = 6'h1b == _myNewVec_59_T_3[5:0] ? myVec_27 : _GEN_388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_390 = 6'h1c == _myNewVec_59_T_3[5:0] ? myVec_28 : _GEN_389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_391 = 6'h1d == _myNewVec_59_T_3[5:0] ? myVec_29 : _GEN_390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_392 = 6'h1e == _myNewVec_59_T_3[5:0] ? myVec_30 : _GEN_391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_393 = 6'h1f == _myNewVec_59_T_3[5:0] ? myVec_31 : _GEN_392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_394 = 6'h20 == _myNewVec_59_T_3[5:0] ? myVec_32 : _GEN_393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_395 = 6'h21 == _myNewVec_59_T_3[5:0] ? myVec_33 : _GEN_394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_396 = 6'h22 == _myNewVec_59_T_3[5:0] ? myVec_34 : _GEN_395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_397 = 6'h23 == _myNewVec_59_T_3[5:0] ? myVec_35 : _GEN_396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_398 = 6'h24 == _myNewVec_59_T_3[5:0] ? myVec_36 : _GEN_397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_399 = 6'h25 == _myNewVec_59_T_3[5:0] ? myVec_37 : _GEN_398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_400 = 6'h26 == _myNewVec_59_T_3[5:0] ? myVec_38 : _GEN_399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_401 = 6'h27 == _myNewVec_59_T_3[5:0] ? myVec_39 : _GEN_400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_402 = 6'h28 == _myNewVec_59_T_3[5:0] ? myVec_40 : _GEN_401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_403 = 6'h29 == _myNewVec_59_T_3[5:0] ? myVec_41 : _GEN_402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_404 = 6'h2a == _myNewVec_59_T_3[5:0] ? myVec_42 : _GEN_403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_405 = 6'h2b == _myNewVec_59_T_3[5:0] ? myVec_43 : _GEN_404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_406 = 6'h2c == _myNewVec_59_T_3[5:0] ? myVec_44 : _GEN_405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_407 = 6'h2d == _myNewVec_59_T_3[5:0] ? myVec_45 : _GEN_406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_408 = 6'h2e == _myNewVec_59_T_3[5:0] ? myVec_46 : _GEN_407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_409 = 6'h2f == _myNewVec_59_T_3[5:0] ? myVec_47 : _GEN_408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_410 = 6'h30 == _myNewVec_59_T_3[5:0] ? myVec_48 : _GEN_409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_411 = 6'h31 == _myNewVec_59_T_3[5:0] ? myVec_49 : _GEN_410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_412 = 6'h32 == _myNewVec_59_T_3[5:0] ? myVec_50 : _GEN_411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_413 = 6'h33 == _myNewVec_59_T_3[5:0] ? myVec_51 : _GEN_412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_414 = 6'h34 == _myNewVec_59_T_3[5:0] ? myVec_52 : _GEN_413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_415 = 6'h35 == _myNewVec_59_T_3[5:0] ? myVec_53 : _GEN_414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_416 = 6'h36 == _myNewVec_59_T_3[5:0] ? myVec_54 : _GEN_415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_417 = 6'h37 == _myNewVec_59_T_3[5:0] ? myVec_55 : _GEN_416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_418 = 6'h38 == _myNewVec_59_T_3[5:0] ? myVec_56 : _GEN_417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_419 = 6'h39 == _myNewVec_59_T_3[5:0] ? myVec_57 : _GEN_418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_420 = 6'h3a == _myNewVec_59_T_3[5:0] ? myVec_58 : _GEN_419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_421 = 6'h3b == _myNewVec_59_T_3[5:0] ? myVec_59 : _GEN_420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_422 = 6'h3c == _myNewVec_59_T_3[5:0] ? myVec_60 : _GEN_421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_423 = 6'h3d == _myNewVec_59_T_3[5:0] ? myVec_61 : _GEN_422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_424 = 6'h3e == _myNewVec_59_T_3[5:0] ? myVec_62 : _GEN_423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_59 = 6'h3f == _myNewVec_59_T_3[5:0] ? myVec_63 : _GEN_424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_58_T_3 = _myNewVec_63_T_1 + 16'h5; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_427 = 6'h1 == _myNewVec_58_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_428 = 6'h2 == _myNewVec_58_T_3[5:0] ? myVec_2 : _GEN_427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_429 = 6'h3 == _myNewVec_58_T_3[5:0] ? myVec_3 : _GEN_428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_430 = 6'h4 == _myNewVec_58_T_3[5:0] ? myVec_4 : _GEN_429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_431 = 6'h5 == _myNewVec_58_T_3[5:0] ? myVec_5 : _GEN_430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_432 = 6'h6 == _myNewVec_58_T_3[5:0] ? myVec_6 : _GEN_431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_433 = 6'h7 == _myNewVec_58_T_3[5:0] ? myVec_7 : _GEN_432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_434 = 6'h8 == _myNewVec_58_T_3[5:0] ? myVec_8 : _GEN_433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_435 = 6'h9 == _myNewVec_58_T_3[5:0] ? myVec_9 : _GEN_434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_436 = 6'ha == _myNewVec_58_T_3[5:0] ? myVec_10 : _GEN_435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_437 = 6'hb == _myNewVec_58_T_3[5:0] ? myVec_11 : _GEN_436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_438 = 6'hc == _myNewVec_58_T_3[5:0] ? myVec_12 : _GEN_437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_439 = 6'hd == _myNewVec_58_T_3[5:0] ? myVec_13 : _GEN_438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_440 = 6'he == _myNewVec_58_T_3[5:0] ? myVec_14 : _GEN_439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_441 = 6'hf == _myNewVec_58_T_3[5:0] ? myVec_15 : _GEN_440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_442 = 6'h10 == _myNewVec_58_T_3[5:0] ? myVec_16 : _GEN_441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_443 = 6'h11 == _myNewVec_58_T_3[5:0] ? myVec_17 : _GEN_442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_444 = 6'h12 == _myNewVec_58_T_3[5:0] ? myVec_18 : _GEN_443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_445 = 6'h13 == _myNewVec_58_T_3[5:0] ? myVec_19 : _GEN_444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_446 = 6'h14 == _myNewVec_58_T_3[5:0] ? myVec_20 : _GEN_445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_447 = 6'h15 == _myNewVec_58_T_3[5:0] ? myVec_21 : _GEN_446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_448 = 6'h16 == _myNewVec_58_T_3[5:0] ? myVec_22 : _GEN_447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_449 = 6'h17 == _myNewVec_58_T_3[5:0] ? myVec_23 : _GEN_448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_450 = 6'h18 == _myNewVec_58_T_3[5:0] ? myVec_24 : _GEN_449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_451 = 6'h19 == _myNewVec_58_T_3[5:0] ? myVec_25 : _GEN_450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_452 = 6'h1a == _myNewVec_58_T_3[5:0] ? myVec_26 : _GEN_451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_453 = 6'h1b == _myNewVec_58_T_3[5:0] ? myVec_27 : _GEN_452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_454 = 6'h1c == _myNewVec_58_T_3[5:0] ? myVec_28 : _GEN_453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_455 = 6'h1d == _myNewVec_58_T_3[5:0] ? myVec_29 : _GEN_454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_456 = 6'h1e == _myNewVec_58_T_3[5:0] ? myVec_30 : _GEN_455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_457 = 6'h1f == _myNewVec_58_T_3[5:0] ? myVec_31 : _GEN_456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_458 = 6'h20 == _myNewVec_58_T_3[5:0] ? myVec_32 : _GEN_457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_459 = 6'h21 == _myNewVec_58_T_3[5:0] ? myVec_33 : _GEN_458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_460 = 6'h22 == _myNewVec_58_T_3[5:0] ? myVec_34 : _GEN_459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_461 = 6'h23 == _myNewVec_58_T_3[5:0] ? myVec_35 : _GEN_460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_462 = 6'h24 == _myNewVec_58_T_3[5:0] ? myVec_36 : _GEN_461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_463 = 6'h25 == _myNewVec_58_T_3[5:0] ? myVec_37 : _GEN_462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_464 = 6'h26 == _myNewVec_58_T_3[5:0] ? myVec_38 : _GEN_463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_465 = 6'h27 == _myNewVec_58_T_3[5:0] ? myVec_39 : _GEN_464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_466 = 6'h28 == _myNewVec_58_T_3[5:0] ? myVec_40 : _GEN_465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_467 = 6'h29 == _myNewVec_58_T_3[5:0] ? myVec_41 : _GEN_466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_468 = 6'h2a == _myNewVec_58_T_3[5:0] ? myVec_42 : _GEN_467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_469 = 6'h2b == _myNewVec_58_T_3[5:0] ? myVec_43 : _GEN_468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_470 = 6'h2c == _myNewVec_58_T_3[5:0] ? myVec_44 : _GEN_469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_471 = 6'h2d == _myNewVec_58_T_3[5:0] ? myVec_45 : _GEN_470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_472 = 6'h2e == _myNewVec_58_T_3[5:0] ? myVec_46 : _GEN_471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_473 = 6'h2f == _myNewVec_58_T_3[5:0] ? myVec_47 : _GEN_472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_474 = 6'h30 == _myNewVec_58_T_3[5:0] ? myVec_48 : _GEN_473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_475 = 6'h31 == _myNewVec_58_T_3[5:0] ? myVec_49 : _GEN_474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_476 = 6'h32 == _myNewVec_58_T_3[5:0] ? myVec_50 : _GEN_475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_477 = 6'h33 == _myNewVec_58_T_3[5:0] ? myVec_51 : _GEN_476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_478 = 6'h34 == _myNewVec_58_T_3[5:0] ? myVec_52 : _GEN_477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_479 = 6'h35 == _myNewVec_58_T_3[5:0] ? myVec_53 : _GEN_478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_480 = 6'h36 == _myNewVec_58_T_3[5:0] ? myVec_54 : _GEN_479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_481 = 6'h37 == _myNewVec_58_T_3[5:0] ? myVec_55 : _GEN_480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_482 = 6'h38 == _myNewVec_58_T_3[5:0] ? myVec_56 : _GEN_481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_483 = 6'h39 == _myNewVec_58_T_3[5:0] ? myVec_57 : _GEN_482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_484 = 6'h3a == _myNewVec_58_T_3[5:0] ? myVec_58 : _GEN_483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_485 = 6'h3b == _myNewVec_58_T_3[5:0] ? myVec_59 : _GEN_484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_486 = 6'h3c == _myNewVec_58_T_3[5:0] ? myVec_60 : _GEN_485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_487 = 6'h3d == _myNewVec_58_T_3[5:0] ? myVec_61 : _GEN_486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_488 = 6'h3e == _myNewVec_58_T_3[5:0] ? myVec_62 : _GEN_487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_58 = 6'h3f == _myNewVec_58_T_3[5:0] ? myVec_63 : _GEN_488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_57_T_3 = _myNewVec_63_T_1 + 16'h6; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_491 = 6'h1 == _myNewVec_57_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_492 = 6'h2 == _myNewVec_57_T_3[5:0] ? myVec_2 : _GEN_491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_493 = 6'h3 == _myNewVec_57_T_3[5:0] ? myVec_3 : _GEN_492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_494 = 6'h4 == _myNewVec_57_T_3[5:0] ? myVec_4 : _GEN_493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_495 = 6'h5 == _myNewVec_57_T_3[5:0] ? myVec_5 : _GEN_494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_496 = 6'h6 == _myNewVec_57_T_3[5:0] ? myVec_6 : _GEN_495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_497 = 6'h7 == _myNewVec_57_T_3[5:0] ? myVec_7 : _GEN_496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_498 = 6'h8 == _myNewVec_57_T_3[5:0] ? myVec_8 : _GEN_497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_499 = 6'h9 == _myNewVec_57_T_3[5:0] ? myVec_9 : _GEN_498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_500 = 6'ha == _myNewVec_57_T_3[5:0] ? myVec_10 : _GEN_499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_501 = 6'hb == _myNewVec_57_T_3[5:0] ? myVec_11 : _GEN_500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_502 = 6'hc == _myNewVec_57_T_3[5:0] ? myVec_12 : _GEN_501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_503 = 6'hd == _myNewVec_57_T_3[5:0] ? myVec_13 : _GEN_502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_504 = 6'he == _myNewVec_57_T_3[5:0] ? myVec_14 : _GEN_503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_505 = 6'hf == _myNewVec_57_T_3[5:0] ? myVec_15 : _GEN_504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_506 = 6'h10 == _myNewVec_57_T_3[5:0] ? myVec_16 : _GEN_505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_507 = 6'h11 == _myNewVec_57_T_3[5:0] ? myVec_17 : _GEN_506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_508 = 6'h12 == _myNewVec_57_T_3[5:0] ? myVec_18 : _GEN_507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_509 = 6'h13 == _myNewVec_57_T_3[5:0] ? myVec_19 : _GEN_508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_510 = 6'h14 == _myNewVec_57_T_3[5:0] ? myVec_20 : _GEN_509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_511 = 6'h15 == _myNewVec_57_T_3[5:0] ? myVec_21 : _GEN_510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_512 = 6'h16 == _myNewVec_57_T_3[5:0] ? myVec_22 : _GEN_511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_513 = 6'h17 == _myNewVec_57_T_3[5:0] ? myVec_23 : _GEN_512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_514 = 6'h18 == _myNewVec_57_T_3[5:0] ? myVec_24 : _GEN_513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_515 = 6'h19 == _myNewVec_57_T_3[5:0] ? myVec_25 : _GEN_514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_516 = 6'h1a == _myNewVec_57_T_3[5:0] ? myVec_26 : _GEN_515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_517 = 6'h1b == _myNewVec_57_T_3[5:0] ? myVec_27 : _GEN_516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_518 = 6'h1c == _myNewVec_57_T_3[5:0] ? myVec_28 : _GEN_517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_519 = 6'h1d == _myNewVec_57_T_3[5:0] ? myVec_29 : _GEN_518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_520 = 6'h1e == _myNewVec_57_T_3[5:0] ? myVec_30 : _GEN_519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_521 = 6'h1f == _myNewVec_57_T_3[5:0] ? myVec_31 : _GEN_520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_522 = 6'h20 == _myNewVec_57_T_3[5:0] ? myVec_32 : _GEN_521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_523 = 6'h21 == _myNewVec_57_T_3[5:0] ? myVec_33 : _GEN_522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_524 = 6'h22 == _myNewVec_57_T_3[5:0] ? myVec_34 : _GEN_523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_525 = 6'h23 == _myNewVec_57_T_3[5:0] ? myVec_35 : _GEN_524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_526 = 6'h24 == _myNewVec_57_T_3[5:0] ? myVec_36 : _GEN_525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_527 = 6'h25 == _myNewVec_57_T_3[5:0] ? myVec_37 : _GEN_526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_528 = 6'h26 == _myNewVec_57_T_3[5:0] ? myVec_38 : _GEN_527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_529 = 6'h27 == _myNewVec_57_T_3[5:0] ? myVec_39 : _GEN_528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_530 = 6'h28 == _myNewVec_57_T_3[5:0] ? myVec_40 : _GEN_529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_531 = 6'h29 == _myNewVec_57_T_3[5:0] ? myVec_41 : _GEN_530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_532 = 6'h2a == _myNewVec_57_T_3[5:0] ? myVec_42 : _GEN_531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_533 = 6'h2b == _myNewVec_57_T_3[5:0] ? myVec_43 : _GEN_532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_534 = 6'h2c == _myNewVec_57_T_3[5:0] ? myVec_44 : _GEN_533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_535 = 6'h2d == _myNewVec_57_T_3[5:0] ? myVec_45 : _GEN_534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_536 = 6'h2e == _myNewVec_57_T_3[5:0] ? myVec_46 : _GEN_535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_537 = 6'h2f == _myNewVec_57_T_3[5:0] ? myVec_47 : _GEN_536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_538 = 6'h30 == _myNewVec_57_T_3[5:0] ? myVec_48 : _GEN_537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_539 = 6'h31 == _myNewVec_57_T_3[5:0] ? myVec_49 : _GEN_538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_540 = 6'h32 == _myNewVec_57_T_3[5:0] ? myVec_50 : _GEN_539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_541 = 6'h33 == _myNewVec_57_T_3[5:0] ? myVec_51 : _GEN_540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_542 = 6'h34 == _myNewVec_57_T_3[5:0] ? myVec_52 : _GEN_541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_543 = 6'h35 == _myNewVec_57_T_3[5:0] ? myVec_53 : _GEN_542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_544 = 6'h36 == _myNewVec_57_T_3[5:0] ? myVec_54 : _GEN_543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_545 = 6'h37 == _myNewVec_57_T_3[5:0] ? myVec_55 : _GEN_544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_546 = 6'h38 == _myNewVec_57_T_3[5:0] ? myVec_56 : _GEN_545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_547 = 6'h39 == _myNewVec_57_T_3[5:0] ? myVec_57 : _GEN_546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_548 = 6'h3a == _myNewVec_57_T_3[5:0] ? myVec_58 : _GEN_547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_549 = 6'h3b == _myNewVec_57_T_3[5:0] ? myVec_59 : _GEN_548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_550 = 6'h3c == _myNewVec_57_T_3[5:0] ? myVec_60 : _GEN_549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_551 = 6'h3d == _myNewVec_57_T_3[5:0] ? myVec_61 : _GEN_550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_552 = 6'h3e == _myNewVec_57_T_3[5:0] ? myVec_62 : _GEN_551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_57 = 6'h3f == _myNewVec_57_T_3[5:0] ? myVec_63 : _GEN_552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_56_T_3 = _myNewVec_63_T_1 + 16'h7; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_555 = 6'h1 == _myNewVec_56_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_556 = 6'h2 == _myNewVec_56_T_3[5:0] ? myVec_2 : _GEN_555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_557 = 6'h3 == _myNewVec_56_T_3[5:0] ? myVec_3 : _GEN_556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_558 = 6'h4 == _myNewVec_56_T_3[5:0] ? myVec_4 : _GEN_557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_559 = 6'h5 == _myNewVec_56_T_3[5:0] ? myVec_5 : _GEN_558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_560 = 6'h6 == _myNewVec_56_T_3[5:0] ? myVec_6 : _GEN_559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_561 = 6'h7 == _myNewVec_56_T_3[5:0] ? myVec_7 : _GEN_560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_562 = 6'h8 == _myNewVec_56_T_3[5:0] ? myVec_8 : _GEN_561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_563 = 6'h9 == _myNewVec_56_T_3[5:0] ? myVec_9 : _GEN_562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_564 = 6'ha == _myNewVec_56_T_3[5:0] ? myVec_10 : _GEN_563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_565 = 6'hb == _myNewVec_56_T_3[5:0] ? myVec_11 : _GEN_564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_566 = 6'hc == _myNewVec_56_T_3[5:0] ? myVec_12 : _GEN_565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_567 = 6'hd == _myNewVec_56_T_3[5:0] ? myVec_13 : _GEN_566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_568 = 6'he == _myNewVec_56_T_3[5:0] ? myVec_14 : _GEN_567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_569 = 6'hf == _myNewVec_56_T_3[5:0] ? myVec_15 : _GEN_568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_570 = 6'h10 == _myNewVec_56_T_3[5:0] ? myVec_16 : _GEN_569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_571 = 6'h11 == _myNewVec_56_T_3[5:0] ? myVec_17 : _GEN_570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_572 = 6'h12 == _myNewVec_56_T_3[5:0] ? myVec_18 : _GEN_571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_573 = 6'h13 == _myNewVec_56_T_3[5:0] ? myVec_19 : _GEN_572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_574 = 6'h14 == _myNewVec_56_T_3[5:0] ? myVec_20 : _GEN_573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_575 = 6'h15 == _myNewVec_56_T_3[5:0] ? myVec_21 : _GEN_574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_576 = 6'h16 == _myNewVec_56_T_3[5:0] ? myVec_22 : _GEN_575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_577 = 6'h17 == _myNewVec_56_T_3[5:0] ? myVec_23 : _GEN_576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_578 = 6'h18 == _myNewVec_56_T_3[5:0] ? myVec_24 : _GEN_577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_579 = 6'h19 == _myNewVec_56_T_3[5:0] ? myVec_25 : _GEN_578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_580 = 6'h1a == _myNewVec_56_T_3[5:0] ? myVec_26 : _GEN_579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_581 = 6'h1b == _myNewVec_56_T_3[5:0] ? myVec_27 : _GEN_580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_582 = 6'h1c == _myNewVec_56_T_3[5:0] ? myVec_28 : _GEN_581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_583 = 6'h1d == _myNewVec_56_T_3[5:0] ? myVec_29 : _GEN_582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_584 = 6'h1e == _myNewVec_56_T_3[5:0] ? myVec_30 : _GEN_583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_585 = 6'h1f == _myNewVec_56_T_3[5:0] ? myVec_31 : _GEN_584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_586 = 6'h20 == _myNewVec_56_T_3[5:0] ? myVec_32 : _GEN_585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_587 = 6'h21 == _myNewVec_56_T_3[5:0] ? myVec_33 : _GEN_586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_588 = 6'h22 == _myNewVec_56_T_3[5:0] ? myVec_34 : _GEN_587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_589 = 6'h23 == _myNewVec_56_T_3[5:0] ? myVec_35 : _GEN_588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_590 = 6'h24 == _myNewVec_56_T_3[5:0] ? myVec_36 : _GEN_589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_591 = 6'h25 == _myNewVec_56_T_3[5:0] ? myVec_37 : _GEN_590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_592 = 6'h26 == _myNewVec_56_T_3[5:0] ? myVec_38 : _GEN_591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_593 = 6'h27 == _myNewVec_56_T_3[5:0] ? myVec_39 : _GEN_592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_594 = 6'h28 == _myNewVec_56_T_3[5:0] ? myVec_40 : _GEN_593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_595 = 6'h29 == _myNewVec_56_T_3[5:0] ? myVec_41 : _GEN_594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_596 = 6'h2a == _myNewVec_56_T_3[5:0] ? myVec_42 : _GEN_595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_597 = 6'h2b == _myNewVec_56_T_3[5:0] ? myVec_43 : _GEN_596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_598 = 6'h2c == _myNewVec_56_T_3[5:0] ? myVec_44 : _GEN_597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_599 = 6'h2d == _myNewVec_56_T_3[5:0] ? myVec_45 : _GEN_598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_600 = 6'h2e == _myNewVec_56_T_3[5:0] ? myVec_46 : _GEN_599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_601 = 6'h2f == _myNewVec_56_T_3[5:0] ? myVec_47 : _GEN_600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_602 = 6'h30 == _myNewVec_56_T_3[5:0] ? myVec_48 : _GEN_601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_603 = 6'h31 == _myNewVec_56_T_3[5:0] ? myVec_49 : _GEN_602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_604 = 6'h32 == _myNewVec_56_T_3[5:0] ? myVec_50 : _GEN_603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_605 = 6'h33 == _myNewVec_56_T_3[5:0] ? myVec_51 : _GEN_604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_606 = 6'h34 == _myNewVec_56_T_3[5:0] ? myVec_52 : _GEN_605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_607 = 6'h35 == _myNewVec_56_T_3[5:0] ? myVec_53 : _GEN_606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_608 = 6'h36 == _myNewVec_56_T_3[5:0] ? myVec_54 : _GEN_607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_609 = 6'h37 == _myNewVec_56_T_3[5:0] ? myVec_55 : _GEN_608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_610 = 6'h38 == _myNewVec_56_T_3[5:0] ? myVec_56 : _GEN_609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_611 = 6'h39 == _myNewVec_56_T_3[5:0] ? myVec_57 : _GEN_610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_612 = 6'h3a == _myNewVec_56_T_3[5:0] ? myVec_58 : _GEN_611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_613 = 6'h3b == _myNewVec_56_T_3[5:0] ? myVec_59 : _GEN_612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_614 = 6'h3c == _myNewVec_56_T_3[5:0] ? myVec_60 : _GEN_613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_615 = 6'h3d == _myNewVec_56_T_3[5:0] ? myVec_61 : _GEN_614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_616 = 6'h3e == _myNewVec_56_T_3[5:0] ? myVec_62 : _GEN_615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_56 = 6'h3f == _myNewVec_56_T_3[5:0] ? myVec_63 : _GEN_616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_55_T_3 = _myNewVec_63_T_1 + 16'h8; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_619 = 6'h1 == _myNewVec_55_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_620 = 6'h2 == _myNewVec_55_T_3[5:0] ? myVec_2 : _GEN_619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_621 = 6'h3 == _myNewVec_55_T_3[5:0] ? myVec_3 : _GEN_620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_622 = 6'h4 == _myNewVec_55_T_3[5:0] ? myVec_4 : _GEN_621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_623 = 6'h5 == _myNewVec_55_T_3[5:0] ? myVec_5 : _GEN_622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_624 = 6'h6 == _myNewVec_55_T_3[5:0] ? myVec_6 : _GEN_623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_625 = 6'h7 == _myNewVec_55_T_3[5:0] ? myVec_7 : _GEN_624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_626 = 6'h8 == _myNewVec_55_T_3[5:0] ? myVec_8 : _GEN_625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_627 = 6'h9 == _myNewVec_55_T_3[5:0] ? myVec_9 : _GEN_626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_628 = 6'ha == _myNewVec_55_T_3[5:0] ? myVec_10 : _GEN_627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_629 = 6'hb == _myNewVec_55_T_3[5:0] ? myVec_11 : _GEN_628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_630 = 6'hc == _myNewVec_55_T_3[5:0] ? myVec_12 : _GEN_629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_631 = 6'hd == _myNewVec_55_T_3[5:0] ? myVec_13 : _GEN_630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_632 = 6'he == _myNewVec_55_T_3[5:0] ? myVec_14 : _GEN_631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_633 = 6'hf == _myNewVec_55_T_3[5:0] ? myVec_15 : _GEN_632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_634 = 6'h10 == _myNewVec_55_T_3[5:0] ? myVec_16 : _GEN_633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_635 = 6'h11 == _myNewVec_55_T_3[5:0] ? myVec_17 : _GEN_634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_636 = 6'h12 == _myNewVec_55_T_3[5:0] ? myVec_18 : _GEN_635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_637 = 6'h13 == _myNewVec_55_T_3[5:0] ? myVec_19 : _GEN_636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_638 = 6'h14 == _myNewVec_55_T_3[5:0] ? myVec_20 : _GEN_637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_639 = 6'h15 == _myNewVec_55_T_3[5:0] ? myVec_21 : _GEN_638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_640 = 6'h16 == _myNewVec_55_T_3[5:0] ? myVec_22 : _GEN_639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_641 = 6'h17 == _myNewVec_55_T_3[5:0] ? myVec_23 : _GEN_640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_642 = 6'h18 == _myNewVec_55_T_3[5:0] ? myVec_24 : _GEN_641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_643 = 6'h19 == _myNewVec_55_T_3[5:0] ? myVec_25 : _GEN_642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_644 = 6'h1a == _myNewVec_55_T_3[5:0] ? myVec_26 : _GEN_643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_645 = 6'h1b == _myNewVec_55_T_3[5:0] ? myVec_27 : _GEN_644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_646 = 6'h1c == _myNewVec_55_T_3[5:0] ? myVec_28 : _GEN_645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_647 = 6'h1d == _myNewVec_55_T_3[5:0] ? myVec_29 : _GEN_646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_648 = 6'h1e == _myNewVec_55_T_3[5:0] ? myVec_30 : _GEN_647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_649 = 6'h1f == _myNewVec_55_T_3[5:0] ? myVec_31 : _GEN_648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_650 = 6'h20 == _myNewVec_55_T_3[5:0] ? myVec_32 : _GEN_649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_651 = 6'h21 == _myNewVec_55_T_3[5:0] ? myVec_33 : _GEN_650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_652 = 6'h22 == _myNewVec_55_T_3[5:0] ? myVec_34 : _GEN_651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_653 = 6'h23 == _myNewVec_55_T_3[5:0] ? myVec_35 : _GEN_652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_654 = 6'h24 == _myNewVec_55_T_3[5:0] ? myVec_36 : _GEN_653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_655 = 6'h25 == _myNewVec_55_T_3[5:0] ? myVec_37 : _GEN_654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_656 = 6'h26 == _myNewVec_55_T_3[5:0] ? myVec_38 : _GEN_655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_657 = 6'h27 == _myNewVec_55_T_3[5:0] ? myVec_39 : _GEN_656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_658 = 6'h28 == _myNewVec_55_T_3[5:0] ? myVec_40 : _GEN_657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_659 = 6'h29 == _myNewVec_55_T_3[5:0] ? myVec_41 : _GEN_658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_660 = 6'h2a == _myNewVec_55_T_3[5:0] ? myVec_42 : _GEN_659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_661 = 6'h2b == _myNewVec_55_T_3[5:0] ? myVec_43 : _GEN_660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_662 = 6'h2c == _myNewVec_55_T_3[5:0] ? myVec_44 : _GEN_661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_663 = 6'h2d == _myNewVec_55_T_3[5:0] ? myVec_45 : _GEN_662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_664 = 6'h2e == _myNewVec_55_T_3[5:0] ? myVec_46 : _GEN_663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_665 = 6'h2f == _myNewVec_55_T_3[5:0] ? myVec_47 : _GEN_664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_666 = 6'h30 == _myNewVec_55_T_3[5:0] ? myVec_48 : _GEN_665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_667 = 6'h31 == _myNewVec_55_T_3[5:0] ? myVec_49 : _GEN_666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_668 = 6'h32 == _myNewVec_55_T_3[5:0] ? myVec_50 : _GEN_667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_669 = 6'h33 == _myNewVec_55_T_3[5:0] ? myVec_51 : _GEN_668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_670 = 6'h34 == _myNewVec_55_T_3[5:0] ? myVec_52 : _GEN_669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_671 = 6'h35 == _myNewVec_55_T_3[5:0] ? myVec_53 : _GEN_670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_672 = 6'h36 == _myNewVec_55_T_3[5:0] ? myVec_54 : _GEN_671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_673 = 6'h37 == _myNewVec_55_T_3[5:0] ? myVec_55 : _GEN_672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_674 = 6'h38 == _myNewVec_55_T_3[5:0] ? myVec_56 : _GEN_673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_675 = 6'h39 == _myNewVec_55_T_3[5:0] ? myVec_57 : _GEN_674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_676 = 6'h3a == _myNewVec_55_T_3[5:0] ? myVec_58 : _GEN_675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_677 = 6'h3b == _myNewVec_55_T_3[5:0] ? myVec_59 : _GEN_676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_678 = 6'h3c == _myNewVec_55_T_3[5:0] ? myVec_60 : _GEN_677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_679 = 6'h3d == _myNewVec_55_T_3[5:0] ? myVec_61 : _GEN_678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_680 = 6'h3e == _myNewVec_55_T_3[5:0] ? myVec_62 : _GEN_679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_55 = 6'h3f == _myNewVec_55_T_3[5:0] ? myVec_63 : _GEN_680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_54_T_3 = _myNewVec_63_T_1 + 16'h9; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_683 = 6'h1 == _myNewVec_54_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_684 = 6'h2 == _myNewVec_54_T_3[5:0] ? myVec_2 : _GEN_683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_685 = 6'h3 == _myNewVec_54_T_3[5:0] ? myVec_3 : _GEN_684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_686 = 6'h4 == _myNewVec_54_T_3[5:0] ? myVec_4 : _GEN_685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_687 = 6'h5 == _myNewVec_54_T_3[5:0] ? myVec_5 : _GEN_686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_688 = 6'h6 == _myNewVec_54_T_3[5:0] ? myVec_6 : _GEN_687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_689 = 6'h7 == _myNewVec_54_T_3[5:0] ? myVec_7 : _GEN_688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_690 = 6'h8 == _myNewVec_54_T_3[5:0] ? myVec_8 : _GEN_689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_691 = 6'h9 == _myNewVec_54_T_3[5:0] ? myVec_9 : _GEN_690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_692 = 6'ha == _myNewVec_54_T_3[5:0] ? myVec_10 : _GEN_691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_693 = 6'hb == _myNewVec_54_T_3[5:0] ? myVec_11 : _GEN_692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_694 = 6'hc == _myNewVec_54_T_3[5:0] ? myVec_12 : _GEN_693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_695 = 6'hd == _myNewVec_54_T_3[5:0] ? myVec_13 : _GEN_694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_696 = 6'he == _myNewVec_54_T_3[5:0] ? myVec_14 : _GEN_695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_697 = 6'hf == _myNewVec_54_T_3[5:0] ? myVec_15 : _GEN_696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_698 = 6'h10 == _myNewVec_54_T_3[5:0] ? myVec_16 : _GEN_697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_699 = 6'h11 == _myNewVec_54_T_3[5:0] ? myVec_17 : _GEN_698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_700 = 6'h12 == _myNewVec_54_T_3[5:0] ? myVec_18 : _GEN_699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_701 = 6'h13 == _myNewVec_54_T_3[5:0] ? myVec_19 : _GEN_700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_702 = 6'h14 == _myNewVec_54_T_3[5:0] ? myVec_20 : _GEN_701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_703 = 6'h15 == _myNewVec_54_T_3[5:0] ? myVec_21 : _GEN_702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_704 = 6'h16 == _myNewVec_54_T_3[5:0] ? myVec_22 : _GEN_703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_705 = 6'h17 == _myNewVec_54_T_3[5:0] ? myVec_23 : _GEN_704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_706 = 6'h18 == _myNewVec_54_T_3[5:0] ? myVec_24 : _GEN_705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_707 = 6'h19 == _myNewVec_54_T_3[5:0] ? myVec_25 : _GEN_706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_708 = 6'h1a == _myNewVec_54_T_3[5:0] ? myVec_26 : _GEN_707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_709 = 6'h1b == _myNewVec_54_T_3[5:0] ? myVec_27 : _GEN_708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_710 = 6'h1c == _myNewVec_54_T_3[5:0] ? myVec_28 : _GEN_709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_711 = 6'h1d == _myNewVec_54_T_3[5:0] ? myVec_29 : _GEN_710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_712 = 6'h1e == _myNewVec_54_T_3[5:0] ? myVec_30 : _GEN_711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_713 = 6'h1f == _myNewVec_54_T_3[5:0] ? myVec_31 : _GEN_712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_714 = 6'h20 == _myNewVec_54_T_3[5:0] ? myVec_32 : _GEN_713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_715 = 6'h21 == _myNewVec_54_T_3[5:0] ? myVec_33 : _GEN_714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_716 = 6'h22 == _myNewVec_54_T_3[5:0] ? myVec_34 : _GEN_715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_717 = 6'h23 == _myNewVec_54_T_3[5:0] ? myVec_35 : _GEN_716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_718 = 6'h24 == _myNewVec_54_T_3[5:0] ? myVec_36 : _GEN_717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_719 = 6'h25 == _myNewVec_54_T_3[5:0] ? myVec_37 : _GEN_718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_720 = 6'h26 == _myNewVec_54_T_3[5:0] ? myVec_38 : _GEN_719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_721 = 6'h27 == _myNewVec_54_T_3[5:0] ? myVec_39 : _GEN_720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_722 = 6'h28 == _myNewVec_54_T_3[5:0] ? myVec_40 : _GEN_721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_723 = 6'h29 == _myNewVec_54_T_3[5:0] ? myVec_41 : _GEN_722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_724 = 6'h2a == _myNewVec_54_T_3[5:0] ? myVec_42 : _GEN_723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_725 = 6'h2b == _myNewVec_54_T_3[5:0] ? myVec_43 : _GEN_724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_726 = 6'h2c == _myNewVec_54_T_3[5:0] ? myVec_44 : _GEN_725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_727 = 6'h2d == _myNewVec_54_T_3[5:0] ? myVec_45 : _GEN_726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_728 = 6'h2e == _myNewVec_54_T_3[5:0] ? myVec_46 : _GEN_727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_729 = 6'h2f == _myNewVec_54_T_3[5:0] ? myVec_47 : _GEN_728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_730 = 6'h30 == _myNewVec_54_T_3[5:0] ? myVec_48 : _GEN_729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_731 = 6'h31 == _myNewVec_54_T_3[5:0] ? myVec_49 : _GEN_730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_732 = 6'h32 == _myNewVec_54_T_3[5:0] ? myVec_50 : _GEN_731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_733 = 6'h33 == _myNewVec_54_T_3[5:0] ? myVec_51 : _GEN_732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_734 = 6'h34 == _myNewVec_54_T_3[5:0] ? myVec_52 : _GEN_733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_735 = 6'h35 == _myNewVec_54_T_3[5:0] ? myVec_53 : _GEN_734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_736 = 6'h36 == _myNewVec_54_T_3[5:0] ? myVec_54 : _GEN_735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_737 = 6'h37 == _myNewVec_54_T_3[5:0] ? myVec_55 : _GEN_736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_738 = 6'h38 == _myNewVec_54_T_3[5:0] ? myVec_56 : _GEN_737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_739 = 6'h39 == _myNewVec_54_T_3[5:0] ? myVec_57 : _GEN_738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_740 = 6'h3a == _myNewVec_54_T_3[5:0] ? myVec_58 : _GEN_739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_741 = 6'h3b == _myNewVec_54_T_3[5:0] ? myVec_59 : _GEN_740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_742 = 6'h3c == _myNewVec_54_T_3[5:0] ? myVec_60 : _GEN_741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_743 = 6'h3d == _myNewVec_54_T_3[5:0] ? myVec_61 : _GEN_742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_744 = 6'h3e == _myNewVec_54_T_3[5:0] ? myVec_62 : _GEN_743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_54 = 6'h3f == _myNewVec_54_T_3[5:0] ? myVec_63 : _GEN_744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_53_T_3 = _myNewVec_63_T_1 + 16'ha; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_747 = 6'h1 == _myNewVec_53_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_748 = 6'h2 == _myNewVec_53_T_3[5:0] ? myVec_2 : _GEN_747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_749 = 6'h3 == _myNewVec_53_T_3[5:0] ? myVec_3 : _GEN_748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_750 = 6'h4 == _myNewVec_53_T_3[5:0] ? myVec_4 : _GEN_749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_751 = 6'h5 == _myNewVec_53_T_3[5:0] ? myVec_5 : _GEN_750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_752 = 6'h6 == _myNewVec_53_T_3[5:0] ? myVec_6 : _GEN_751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_753 = 6'h7 == _myNewVec_53_T_3[5:0] ? myVec_7 : _GEN_752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_754 = 6'h8 == _myNewVec_53_T_3[5:0] ? myVec_8 : _GEN_753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_755 = 6'h9 == _myNewVec_53_T_3[5:0] ? myVec_9 : _GEN_754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_756 = 6'ha == _myNewVec_53_T_3[5:0] ? myVec_10 : _GEN_755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_757 = 6'hb == _myNewVec_53_T_3[5:0] ? myVec_11 : _GEN_756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_758 = 6'hc == _myNewVec_53_T_3[5:0] ? myVec_12 : _GEN_757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_759 = 6'hd == _myNewVec_53_T_3[5:0] ? myVec_13 : _GEN_758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_760 = 6'he == _myNewVec_53_T_3[5:0] ? myVec_14 : _GEN_759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_761 = 6'hf == _myNewVec_53_T_3[5:0] ? myVec_15 : _GEN_760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_762 = 6'h10 == _myNewVec_53_T_3[5:0] ? myVec_16 : _GEN_761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_763 = 6'h11 == _myNewVec_53_T_3[5:0] ? myVec_17 : _GEN_762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_764 = 6'h12 == _myNewVec_53_T_3[5:0] ? myVec_18 : _GEN_763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_765 = 6'h13 == _myNewVec_53_T_3[5:0] ? myVec_19 : _GEN_764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_766 = 6'h14 == _myNewVec_53_T_3[5:0] ? myVec_20 : _GEN_765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_767 = 6'h15 == _myNewVec_53_T_3[5:0] ? myVec_21 : _GEN_766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_768 = 6'h16 == _myNewVec_53_T_3[5:0] ? myVec_22 : _GEN_767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_769 = 6'h17 == _myNewVec_53_T_3[5:0] ? myVec_23 : _GEN_768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_770 = 6'h18 == _myNewVec_53_T_3[5:0] ? myVec_24 : _GEN_769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_771 = 6'h19 == _myNewVec_53_T_3[5:0] ? myVec_25 : _GEN_770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_772 = 6'h1a == _myNewVec_53_T_3[5:0] ? myVec_26 : _GEN_771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_773 = 6'h1b == _myNewVec_53_T_3[5:0] ? myVec_27 : _GEN_772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_774 = 6'h1c == _myNewVec_53_T_3[5:0] ? myVec_28 : _GEN_773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_775 = 6'h1d == _myNewVec_53_T_3[5:0] ? myVec_29 : _GEN_774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_776 = 6'h1e == _myNewVec_53_T_3[5:0] ? myVec_30 : _GEN_775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_777 = 6'h1f == _myNewVec_53_T_3[5:0] ? myVec_31 : _GEN_776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_778 = 6'h20 == _myNewVec_53_T_3[5:0] ? myVec_32 : _GEN_777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_779 = 6'h21 == _myNewVec_53_T_3[5:0] ? myVec_33 : _GEN_778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_780 = 6'h22 == _myNewVec_53_T_3[5:0] ? myVec_34 : _GEN_779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_781 = 6'h23 == _myNewVec_53_T_3[5:0] ? myVec_35 : _GEN_780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_782 = 6'h24 == _myNewVec_53_T_3[5:0] ? myVec_36 : _GEN_781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_783 = 6'h25 == _myNewVec_53_T_3[5:0] ? myVec_37 : _GEN_782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_784 = 6'h26 == _myNewVec_53_T_3[5:0] ? myVec_38 : _GEN_783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_785 = 6'h27 == _myNewVec_53_T_3[5:0] ? myVec_39 : _GEN_784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_786 = 6'h28 == _myNewVec_53_T_3[5:0] ? myVec_40 : _GEN_785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_787 = 6'h29 == _myNewVec_53_T_3[5:0] ? myVec_41 : _GEN_786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_788 = 6'h2a == _myNewVec_53_T_3[5:0] ? myVec_42 : _GEN_787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_789 = 6'h2b == _myNewVec_53_T_3[5:0] ? myVec_43 : _GEN_788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_790 = 6'h2c == _myNewVec_53_T_3[5:0] ? myVec_44 : _GEN_789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_791 = 6'h2d == _myNewVec_53_T_3[5:0] ? myVec_45 : _GEN_790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_792 = 6'h2e == _myNewVec_53_T_3[5:0] ? myVec_46 : _GEN_791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_793 = 6'h2f == _myNewVec_53_T_3[5:0] ? myVec_47 : _GEN_792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_794 = 6'h30 == _myNewVec_53_T_3[5:0] ? myVec_48 : _GEN_793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_795 = 6'h31 == _myNewVec_53_T_3[5:0] ? myVec_49 : _GEN_794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_796 = 6'h32 == _myNewVec_53_T_3[5:0] ? myVec_50 : _GEN_795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_797 = 6'h33 == _myNewVec_53_T_3[5:0] ? myVec_51 : _GEN_796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_798 = 6'h34 == _myNewVec_53_T_3[5:0] ? myVec_52 : _GEN_797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_799 = 6'h35 == _myNewVec_53_T_3[5:0] ? myVec_53 : _GEN_798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_800 = 6'h36 == _myNewVec_53_T_3[5:0] ? myVec_54 : _GEN_799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_801 = 6'h37 == _myNewVec_53_T_3[5:0] ? myVec_55 : _GEN_800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_802 = 6'h38 == _myNewVec_53_T_3[5:0] ? myVec_56 : _GEN_801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_803 = 6'h39 == _myNewVec_53_T_3[5:0] ? myVec_57 : _GEN_802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_804 = 6'h3a == _myNewVec_53_T_3[5:0] ? myVec_58 : _GEN_803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_805 = 6'h3b == _myNewVec_53_T_3[5:0] ? myVec_59 : _GEN_804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_806 = 6'h3c == _myNewVec_53_T_3[5:0] ? myVec_60 : _GEN_805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_807 = 6'h3d == _myNewVec_53_T_3[5:0] ? myVec_61 : _GEN_806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_808 = 6'h3e == _myNewVec_53_T_3[5:0] ? myVec_62 : _GEN_807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_53 = 6'h3f == _myNewVec_53_T_3[5:0] ? myVec_63 : _GEN_808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_52_T_3 = _myNewVec_63_T_1 + 16'hb; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_811 = 6'h1 == _myNewVec_52_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_812 = 6'h2 == _myNewVec_52_T_3[5:0] ? myVec_2 : _GEN_811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_813 = 6'h3 == _myNewVec_52_T_3[5:0] ? myVec_3 : _GEN_812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_814 = 6'h4 == _myNewVec_52_T_3[5:0] ? myVec_4 : _GEN_813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_815 = 6'h5 == _myNewVec_52_T_3[5:0] ? myVec_5 : _GEN_814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_816 = 6'h6 == _myNewVec_52_T_3[5:0] ? myVec_6 : _GEN_815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_817 = 6'h7 == _myNewVec_52_T_3[5:0] ? myVec_7 : _GEN_816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_818 = 6'h8 == _myNewVec_52_T_3[5:0] ? myVec_8 : _GEN_817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_819 = 6'h9 == _myNewVec_52_T_3[5:0] ? myVec_9 : _GEN_818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_820 = 6'ha == _myNewVec_52_T_3[5:0] ? myVec_10 : _GEN_819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_821 = 6'hb == _myNewVec_52_T_3[5:0] ? myVec_11 : _GEN_820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_822 = 6'hc == _myNewVec_52_T_3[5:0] ? myVec_12 : _GEN_821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_823 = 6'hd == _myNewVec_52_T_3[5:0] ? myVec_13 : _GEN_822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_824 = 6'he == _myNewVec_52_T_3[5:0] ? myVec_14 : _GEN_823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_825 = 6'hf == _myNewVec_52_T_3[5:0] ? myVec_15 : _GEN_824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_826 = 6'h10 == _myNewVec_52_T_3[5:0] ? myVec_16 : _GEN_825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_827 = 6'h11 == _myNewVec_52_T_3[5:0] ? myVec_17 : _GEN_826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_828 = 6'h12 == _myNewVec_52_T_3[5:0] ? myVec_18 : _GEN_827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_829 = 6'h13 == _myNewVec_52_T_3[5:0] ? myVec_19 : _GEN_828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_830 = 6'h14 == _myNewVec_52_T_3[5:0] ? myVec_20 : _GEN_829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_831 = 6'h15 == _myNewVec_52_T_3[5:0] ? myVec_21 : _GEN_830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_832 = 6'h16 == _myNewVec_52_T_3[5:0] ? myVec_22 : _GEN_831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_833 = 6'h17 == _myNewVec_52_T_3[5:0] ? myVec_23 : _GEN_832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_834 = 6'h18 == _myNewVec_52_T_3[5:0] ? myVec_24 : _GEN_833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_835 = 6'h19 == _myNewVec_52_T_3[5:0] ? myVec_25 : _GEN_834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_836 = 6'h1a == _myNewVec_52_T_3[5:0] ? myVec_26 : _GEN_835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_837 = 6'h1b == _myNewVec_52_T_3[5:0] ? myVec_27 : _GEN_836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_838 = 6'h1c == _myNewVec_52_T_3[5:0] ? myVec_28 : _GEN_837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_839 = 6'h1d == _myNewVec_52_T_3[5:0] ? myVec_29 : _GEN_838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_840 = 6'h1e == _myNewVec_52_T_3[5:0] ? myVec_30 : _GEN_839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_841 = 6'h1f == _myNewVec_52_T_3[5:0] ? myVec_31 : _GEN_840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_842 = 6'h20 == _myNewVec_52_T_3[5:0] ? myVec_32 : _GEN_841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_843 = 6'h21 == _myNewVec_52_T_3[5:0] ? myVec_33 : _GEN_842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_844 = 6'h22 == _myNewVec_52_T_3[5:0] ? myVec_34 : _GEN_843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_845 = 6'h23 == _myNewVec_52_T_3[5:0] ? myVec_35 : _GEN_844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_846 = 6'h24 == _myNewVec_52_T_3[5:0] ? myVec_36 : _GEN_845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_847 = 6'h25 == _myNewVec_52_T_3[5:0] ? myVec_37 : _GEN_846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_848 = 6'h26 == _myNewVec_52_T_3[5:0] ? myVec_38 : _GEN_847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_849 = 6'h27 == _myNewVec_52_T_3[5:0] ? myVec_39 : _GEN_848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_850 = 6'h28 == _myNewVec_52_T_3[5:0] ? myVec_40 : _GEN_849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_851 = 6'h29 == _myNewVec_52_T_3[5:0] ? myVec_41 : _GEN_850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_852 = 6'h2a == _myNewVec_52_T_3[5:0] ? myVec_42 : _GEN_851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_853 = 6'h2b == _myNewVec_52_T_3[5:0] ? myVec_43 : _GEN_852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_854 = 6'h2c == _myNewVec_52_T_3[5:0] ? myVec_44 : _GEN_853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_855 = 6'h2d == _myNewVec_52_T_3[5:0] ? myVec_45 : _GEN_854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_856 = 6'h2e == _myNewVec_52_T_3[5:0] ? myVec_46 : _GEN_855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_857 = 6'h2f == _myNewVec_52_T_3[5:0] ? myVec_47 : _GEN_856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_858 = 6'h30 == _myNewVec_52_T_3[5:0] ? myVec_48 : _GEN_857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_859 = 6'h31 == _myNewVec_52_T_3[5:0] ? myVec_49 : _GEN_858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_860 = 6'h32 == _myNewVec_52_T_3[5:0] ? myVec_50 : _GEN_859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_861 = 6'h33 == _myNewVec_52_T_3[5:0] ? myVec_51 : _GEN_860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_862 = 6'h34 == _myNewVec_52_T_3[5:0] ? myVec_52 : _GEN_861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_863 = 6'h35 == _myNewVec_52_T_3[5:0] ? myVec_53 : _GEN_862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_864 = 6'h36 == _myNewVec_52_T_3[5:0] ? myVec_54 : _GEN_863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_865 = 6'h37 == _myNewVec_52_T_3[5:0] ? myVec_55 : _GEN_864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_866 = 6'h38 == _myNewVec_52_T_3[5:0] ? myVec_56 : _GEN_865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_867 = 6'h39 == _myNewVec_52_T_3[5:0] ? myVec_57 : _GEN_866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_868 = 6'h3a == _myNewVec_52_T_3[5:0] ? myVec_58 : _GEN_867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_869 = 6'h3b == _myNewVec_52_T_3[5:0] ? myVec_59 : _GEN_868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_870 = 6'h3c == _myNewVec_52_T_3[5:0] ? myVec_60 : _GEN_869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_871 = 6'h3d == _myNewVec_52_T_3[5:0] ? myVec_61 : _GEN_870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_872 = 6'h3e == _myNewVec_52_T_3[5:0] ? myVec_62 : _GEN_871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_52 = 6'h3f == _myNewVec_52_T_3[5:0] ? myVec_63 : _GEN_872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_51_T_3 = _myNewVec_63_T_1 + 16'hc; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_875 = 6'h1 == _myNewVec_51_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_876 = 6'h2 == _myNewVec_51_T_3[5:0] ? myVec_2 : _GEN_875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_877 = 6'h3 == _myNewVec_51_T_3[5:0] ? myVec_3 : _GEN_876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_878 = 6'h4 == _myNewVec_51_T_3[5:0] ? myVec_4 : _GEN_877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_879 = 6'h5 == _myNewVec_51_T_3[5:0] ? myVec_5 : _GEN_878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_880 = 6'h6 == _myNewVec_51_T_3[5:0] ? myVec_6 : _GEN_879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_881 = 6'h7 == _myNewVec_51_T_3[5:0] ? myVec_7 : _GEN_880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_882 = 6'h8 == _myNewVec_51_T_3[5:0] ? myVec_8 : _GEN_881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_883 = 6'h9 == _myNewVec_51_T_3[5:0] ? myVec_9 : _GEN_882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_884 = 6'ha == _myNewVec_51_T_3[5:0] ? myVec_10 : _GEN_883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_885 = 6'hb == _myNewVec_51_T_3[5:0] ? myVec_11 : _GEN_884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_886 = 6'hc == _myNewVec_51_T_3[5:0] ? myVec_12 : _GEN_885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_887 = 6'hd == _myNewVec_51_T_3[5:0] ? myVec_13 : _GEN_886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_888 = 6'he == _myNewVec_51_T_3[5:0] ? myVec_14 : _GEN_887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_889 = 6'hf == _myNewVec_51_T_3[5:0] ? myVec_15 : _GEN_888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_890 = 6'h10 == _myNewVec_51_T_3[5:0] ? myVec_16 : _GEN_889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_891 = 6'h11 == _myNewVec_51_T_3[5:0] ? myVec_17 : _GEN_890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_892 = 6'h12 == _myNewVec_51_T_3[5:0] ? myVec_18 : _GEN_891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_893 = 6'h13 == _myNewVec_51_T_3[5:0] ? myVec_19 : _GEN_892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_894 = 6'h14 == _myNewVec_51_T_3[5:0] ? myVec_20 : _GEN_893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_895 = 6'h15 == _myNewVec_51_T_3[5:0] ? myVec_21 : _GEN_894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_896 = 6'h16 == _myNewVec_51_T_3[5:0] ? myVec_22 : _GEN_895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_897 = 6'h17 == _myNewVec_51_T_3[5:0] ? myVec_23 : _GEN_896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_898 = 6'h18 == _myNewVec_51_T_3[5:0] ? myVec_24 : _GEN_897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_899 = 6'h19 == _myNewVec_51_T_3[5:0] ? myVec_25 : _GEN_898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_900 = 6'h1a == _myNewVec_51_T_3[5:0] ? myVec_26 : _GEN_899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_901 = 6'h1b == _myNewVec_51_T_3[5:0] ? myVec_27 : _GEN_900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_902 = 6'h1c == _myNewVec_51_T_3[5:0] ? myVec_28 : _GEN_901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_903 = 6'h1d == _myNewVec_51_T_3[5:0] ? myVec_29 : _GEN_902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_904 = 6'h1e == _myNewVec_51_T_3[5:0] ? myVec_30 : _GEN_903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_905 = 6'h1f == _myNewVec_51_T_3[5:0] ? myVec_31 : _GEN_904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_906 = 6'h20 == _myNewVec_51_T_3[5:0] ? myVec_32 : _GEN_905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_907 = 6'h21 == _myNewVec_51_T_3[5:0] ? myVec_33 : _GEN_906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_908 = 6'h22 == _myNewVec_51_T_3[5:0] ? myVec_34 : _GEN_907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_909 = 6'h23 == _myNewVec_51_T_3[5:0] ? myVec_35 : _GEN_908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_910 = 6'h24 == _myNewVec_51_T_3[5:0] ? myVec_36 : _GEN_909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_911 = 6'h25 == _myNewVec_51_T_3[5:0] ? myVec_37 : _GEN_910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_912 = 6'h26 == _myNewVec_51_T_3[5:0] ? myVec_38 : _GEN_911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_913 = 6'h27 == _myNewVec_51_T_3[5:0] ? myVec_39 : _GEN_912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_914 = 6'h28 == _myNewVec_51_T_3[5:0] ? myVec_40 : _GEN_913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_915 = 6'h29 == _myNewVec_51_T_3[5:0] ? myVec_41 : _GEN_914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_916 = 6'h2a == _myNewVec_51_T_3[5:0] ? myVec_42 : _GEN_915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_917 = 6'h2b == _myNewVec_51_T_3[5:0] ? myVec_43 : _GEN_916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_918 = 6'h2c == _myNewVec_51_T_3[5:0] ? myVec_44 : _GEN_917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_919 = 6'h2d == _myNewVec_51_T_3[5:0] ? myVec_45 : _GEN_918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_920 = 6'h2e == _myNewVec_51_T_3[5:0] ? myVec_46 : _GEN_919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_921 = 6'h2f == _myNewVec_51_T_3[5:0] ? myVec_47 : _GEN_920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_922 = 6'h30 == _myNewVec_51_T_3[5:0] ? myVec_48 : _GEN_921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_923 = 6'h31 == _myNewVec_51_T_3[5:0] ? myVec_49 : _GEN_922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_924 = 6'h32 == _myNewVec_51_T_3[5:0] ? myVec_50 : _GEN_923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_925 = 6'h33 == _myNewVec_51_T_3[5:0] ? myVec_51 : _GEN_924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_926 = 6'h34 == _myNewVec_51_T_3[5:0] ? myVec_52 : _GEN_925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_927 = 6'h35 == _myNewVec_51_T_3[5:0] ? myVec_53 : _GEN_926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_928 = 6'h36 == _myNewVec_51_T_3[5:0] ? myVec_54 : _GEN_927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_929 = 6'h37 == _myNewVec_51_T_3[5:0] ? myVec_55 : _GEN_928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_930 = 6'h38 == _myNewVec_51_T_3[5:0] ? myVec_56 : _GEN_929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_931 = 6'h39 == _myNewVec_51_T_3[5:0] ? myVec_57 : _GEN_930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_932 = 6'h3a == _myNewVec_51_T_3[5:0] ? myVec_58 : _GEN_931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_933 = 6'h3b == _myNewVec_51_T_3[5:0] ? myVec_59 : _GEN_932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_934 = 6'h3c == _myNewVec_51_T_3[5:0] ? myVec_60 : _GEN_933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_935 = 6'h3d == _myNewVec_51_T_3[5:0] ? myVec_61 : _GEN_934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_936 = 6'h3e == _myNewVec_51_T_3[5:0] ? myVec_62 : _GEN_935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_51 = 6'h3f == _myNewVec_51_T_3[5:0] ? myVec_63 : _GEN_936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_50_T_3 = _myNewVec_63_T_1 + 16'hd; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_939 = 6'h1 == _myNewVec_50_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_940 = 6'h2 == _myNewVec_50_T_3[5:0] ? myVec_2 : _GEN_939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_941 = 6'h3 == _myNewVec_50_T_3[5:0] ? myVec_3 : _GEN_940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_942 = 6'h4 == _myNewVec_50_T_3[5:0] ? myVec_4 : _GEN_941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_943 = 6'h5 == _myNewVec_50_T_3[5:0] ? myVec_5 : _GEN_942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_944 = 6'h6 == _myNewVec_50_T_3[5:0] ? myVec_6 : _GEN_943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_945 = 6'h7 == _myNewVec_50_T_3[5:0] ? myVec_7 : _GEN_944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_946 = 6'h8 == _myNewVec_50_T_3[5:0] ? myVec_8 : _GEN_945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_947 = 6'h9 == _myNewVec_50_T_3[5:0] ? myVec_9 : _GEN_946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_948 = 6'ha == _myNewVec_50_T_3[5:0] ? myVec_10 : _GEN_947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_949 = 6'hb == _myNewVec_50_T_3[5:0] ? myVec_11 : _GEN_948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_950 = 6'hc == _myNewVec_50_T_3[5:0] ? myVec_12 : _GEN_949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_951 = 6'hd == _myNewVec_50_T_3[5:0] ? myVec_13 : _GEN_950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_952 = 6'he == _myNewVec_50_T_3[5:0] ? myVec_14 : _GEN_951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_953 = 6'hf == _myNewVec_50_T_3[5:0] ? myVec_15 : _GEN_952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_954 = 6'h10 == _myNewVec_50_T_3[5:0] ? myVec_16 : _GEN_953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_955 = 6'h11 == _myNewVec_50_T_3[5:0] ? myVec_17 : _GEN_954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_956 = 6'h12 == _myNewVec_50_T_3[5:0] ? myVec_18 : _GEN_955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_957 = 6'h13 == _myNewVec_50_T_3[5:0] ? myVec_19 : _GEN_956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_958 = 6'h14 == _myNewVec_50_T_3[5:0] ? myVec_20 : _GEN_957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_959 = 6'h15 == _myNewVec_50_T_3[5:0] ? myVec_21 : _GEN_958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_960 = 6'h16 == _myNewVec_50_T_3[5:0] ? myVec_22 : _GEN_959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_961 = 6'h17 == _myNewVec_50_T_3[5:0] ? myVec_23 : _GEN_960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_962 = 6'h18 == _myNewVec_50_T_3[5:0] ? myVec_24 : _GEN_961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_963 = 6'h19 == _myNewVec_50_T_3[5:0] ? myVec_25 : _GEN_962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_964 = 6'h1a == _myNewVec_50_T_3[5:0] ? myVec_26 : _GEN_963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_965 = 6'h1b == _myNewVec_50_T_3[5:0] ? myVec_27 : _GEN_964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_966 = 6'h1c == _myNewVec_50_T_3[5:0] ? myVec_28 : _GEN_965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_967 = 6'h1d == _myNewVec_50_T_3[5:0] ? myVec_29 : _GEN_966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_968 = 6'h1e == _myNewVec_50_T_3[5:0] ? myVec_30 : _GEN_967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_969 = 6'h1f == _myNewVec_50_T_3[5:0] ? myVec_31 : _GEN_968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_970 = 6'h20 == _myNewVec_50_T_3[5:0] ? myVec_32 : _GEN_969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_971 = 6'h21 == _myNewVec_50_T_3[5:0] ? myVec_33 : _GEN_970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_972 = 6'h22 == _myNewVec_50_T_3[5:0] ? myVec_34 : _GEN_971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_973 = 6'h23 == _myNewVec_50_T_3[5:0] ? myVec_35 : _GEN_972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_974 = 6'h24 == _myNewVec_50_T_3[5:0] ? myVec_36 : _GEN_973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_975 = 6'h25 == _myNewVec_50_T_3[5:0] ? myVec_37 : _GEN_974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_976 = 6'h26 == _myNewVec_50_T_3[5:0] ? myVec_38 : _GEN_975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_977 = 6'h27 == _myNewVec_50_T_3[5:0] ? myVec_39 : _GEN_976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_978 = 6'h28 == _myNewVec_50_T_3[5:0] ? myVec_40 : _GEN_977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_979 = 6'h29 == _myNewVec_50_T_3[5:0] ? myVec_41 : _GEN_978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_980 = 6'h2a == _myNewVec_50_T_3[5:0] ? myVec_42 : _GEN_979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_981 = 6'h2b == _myNewVec_50_T_3[5:0] ? myVec_43 : _GEN_980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_982 = 6'h2c == _myNewVec_50_T_3[5:0] ? myVec_44 : _GEN_981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_983 = 6'h2d == _myNewVec_50_T_3[5:0] ? myVec_45 : _GEN_982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_984 = 6'h2e == _myNewVec_50_T_3[5:0] ? myVec_46 : _GEN_983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_985 = 6'h2f == _myNewVec_50_T_3[5:0] ? myVec_47 : _GEN_984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_986 = 6'h30 == _myNewVec_50_T_3[5:0] ? myVec_48 : _GEN_985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_987 = 6'h31 == _myNewVec_50_T_3[5:0] ? myVec_49 : _GEN_986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_988 = 6'h32 == _myNewVec_50_T_3[5:0] ? myVec_50 : _GEN_987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_989 = 6'h33 == _myNewVec_50_T_3[5:0] ? myVec_51 : _GEN_988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_990 = 6'h34 == _myNewVec_50_T_3[5:0] ? myVec_52 : _GEN_989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_991 = 6'h35 == _myNewVec_50_T_3[5:0] ? myVec_53 : _GEN_990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_992 = 6'h36 == _myNewVec_50_T_3[5:0] ? myVec_54 : _GEN_991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_993 = 6'h37 == _myNewVec_50_T_3[5:0] ? myVec_55 : _GEN_992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_994 = 6'h38 == _myNewVec_50_T_3[5:0] ? myVec_56 : _GEN_993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_995 = 6'h39 == _myNewVec_50_T_3[5:0] ? myVec_57 : _GEN_994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_996 = 6'h3a == _myNewVec_50_T_3[5:0] ? myVec_58 : _GEN_995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_997 = 6'h3b == _myNewVec_50_T_3[5:0] ? myVec_59 : _GEN_996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_998 = 6'h3c == _myNewVec_50_T_3[5:0] ? myVec_60 : _GEN_997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_999 = 6'h3d == _myNewVec_50_T_3[5:0] ? myVec_61 : _GEN_998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1000 = 6'h3e == _myNewVec_50_T_3[5:0] ? myVec_62 : _GEN_999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_50 = 6'h3f == _myNewVec_50_T_3[5:0] ? myVec_63 : _GEN_1000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_49_T_3 = _myNewVec_63_T_1 + 16'he; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1003 = 6'h1 == _myNewVec_49_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1004 = 6'h2 == _myNewVec_49_T_3[5:0] ? myVec_2 : _GEN_1003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1005 = 6'h3 == _myNewVec_49_T_3[5:0] ? myVec_3 : _GEN_1004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1006 = 6'h4 == _myNewVec_49_T_3[5:0] ? myVec_4 : _GEN_1005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1007 = 6'h5 == _myNewVec_49_T_3[5:0] ? myVec_5 : _GEN_1006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1008 = 6'h6 == _myNewVec_49_T_3[5:0] ? myVec_6 : _GEN_1007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1009 = 6'h7 == _myNewVec_49_T_3[5:0] ? myVec_7 : _GEN_1008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1010 = 6'h8 == _myNewVec_49_T_3[5:0] ? myVec_8 : _GEN_1009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1011 = 6'h9 == _myNewVec_49_T_3[5:0] ? myVec_9 : _GEN_1010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1012 = 6'ha == _myNewVec_49_T_3[5:0] ? myVec_10 : _GEN_1011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1013 = 6'hb == _myNewVec_49_T_3[5:0] ? myVec_11 : _GEN_1012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1014 = 6'hc == _myNewVec_49_T_3[5:0] ? myVec_12 : _GEN_1013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1015 = 6'hd == _myNewVec_49_T_3[5:0] ? myVec_13 : _GEN_1014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1016 = 6'he == _myNewVec_49_T_3[5:0] ? myVec_14 : _GEN_1015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1017 = 6'hf == _myNewVec_49_T_3[5:0] ? myVec_15 : _GEN_1016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1018 = 6'h10 == _myNewVec_49_T_3[5:0] ? myVec_16 : _GEN_1017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1019 = 6'h11 == _myNewVec_49_T_3[5:0] ? myVec_17 : _GEN_1018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1020 = 6'h12 == _myNewVec_49_T_3[5:0] ? myVec_18 : _GEN_1019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1021 = 6'h13 == _myNewVec_49_T_3[5:0] ? myVec_19 : _GEN_1020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1022 = 6'h14 == _myNewVec_49_T_3[5:0] ? myVec_20 : _GEN_1021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1023 = 6'h15 == _myNewVec_49_T_3[5:0] ? myVec_21 : _GEN_1022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1024 = 6'h16 == _myNewVec_49_T_3[5:0] ? myVec_22 : _GEN_1023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1025 = 6'h17 == _myNewVec_49_T_3[5:0] ? myVec_23 : _GEN_1024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1026 = 6'h18 == _myNewVec_49_T_3[5:0] ? myVec_24 : _GEN_1025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1027 = 6'h19 == _myNewVec_49_T_3[5:0] ? myVec_25 : _GEN_1026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1028 = 6'h1a == _myNewVec_49_T_3[5:0] ? myVec_26 : _GEN_1027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1029 = 6'h1b == _myNewVec_49_T_3[5:0] ? myVec_27 : _GEN_1028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1030 = 6'h1c == _myNewVec_49_T_3[5:0] ? myVec_28 : _GEN_1029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1031 = 6'h1d == _myNewVec_49_T_3[5:0] ? myVec_29 : _GEN_1030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1032 = 6'h1e == _myNewVec_49_T_3[5:0] ? myVec_30 : _GEN_1031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1033 = 6'h1f == _myNewVec_49_T_3[5:0] ? myVec_31 : _GEN_1032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1034 = 6'h20 == _myNewVec_49_T_3[5:0] ? myVec_32 : _GEN_1033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1035 = 6'h21 == _myNewVec_49_T_3[5:0] ? myVec_33 : _GEN_1034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1036 = 6'h22 == _myNewVec_49_T_3[5:0] ? myVec_34 : _GEN_1035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1037 = 6'h23 == _myNewVec_49_T_3[5:0] ? myVec_35 : _GEN_1036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1038 = 6'h24 == _myNewVec_49_T_3[5:0] ? myVec_36 : _GEN_1037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1039 = 6'h25 == _myNewVec_49_T_3[5:0] ? myVec_37 : _GEN_1038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1040 = 6'h26 == _myNewVec_49_T_3[5:0] ? myVec_38 : _GEN_1039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1041 = 6'h27 == _myNewVec_49_T_3[5:0] ? myVec_39 : _GEN_1040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1042 = 6'h28 == _myNewVec_49_T_3[5:0] ? myVec_40 : _GEN_1041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1043 = 6'h29 == _myNewVec_49_T_3[5:0] ? myVec_41 : _GEN_1042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1044 = 6'h2a == _myNewVec_49_T_3[5:0] ? myVec_42 : _GEN_1043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1045 = 6'h2b == _myNewVec_49_T_3[5:0] ? myVec_43 : _GEN_1044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1046 = 6'h2c == _myNewVec_49_T_3[5:0] ? myVec_44 : _GEN_1045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1047 = 6'h2d == _myNewVec_49_T_3[5:0] ? myVec_45 : _GEN_1046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1048 = 6'h2e == _myNewVec_49_T_3[5:0] ? myVec_46 : _GEN_1047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1049 = 6'h2f == _myNewVec_49_T_3[5:0] ? myVec_47 : _GEN_1048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1050 = 6'h30 == _myNewVec_49_T_3[5:0] ? myVec_48 : _GEN_1049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1051 = 6'h31 == _myNewVec_49_T_3[5:0] ? myVec_49 : _GEN_1050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1052 = 6'h32 == _myNewVec_49_T_3[5:0] ? myVec_50 : _GEN_1051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1053 = 6'h33 == _myNewVec_49_T_3[5:0] ? myVec_51 : _GEN_1052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1054 = 6'h34 == _myNewVec_49_T_3[5:0] ? myVec_52 : _GEN_1053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1055 = 6'h35 == _myNewVec_49_T_3[5:0] ? myVec_53 : _GEN_1054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1056 = 6'h36 == _myNewVec_49_T_3[5:0] ? myVec_54 : _GEN_1055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1057 = 6'h37 == _myNewVec_49_T_3[5:0] ? myVec_55 : _GEN_1056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1058 = 6'h38 == _myNewVec_49_T_3[5:0] ? myVec_56 : _GEN_1057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1059 = 6'h39 == _myNewVec_49_T_3[5:0] ? myVec_57 : _GEN_1058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1060 = 6'h3a == _myNewVec_49_T_3[5:0] ? myVec_58 : _GEN_1059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1061 = 6'h3b == _myNewVec_49_T_3[5:0] ? myVec_59 : _GEN_1060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1062 = 6'h3c == _myNewVec_49_T_3[5:0] ? myVec_60 : _GEN_1061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1063 = 6'h3d == _myNewVec_49_T_3[5:0] ? myVec_61 : _GEN_1062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1064 = 6'h3e == _myNewVec_49_T_3[5:0] ? myVec_62 : _GEN_1063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_49 = 6'h3f == _myNewVec_49_T_3[5:0] ? myVec_63 : _GEN_1064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_48_T_3 = _myNewVec_63_T_1 + 16'hf; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1067 = 6'h1 == _myNewVec_48_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1068 = 6'h2 == _myNewVec_48_T_3[5:0] ? myVec_2 : _GEN_1067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1069 = 6'h3 == _myNewVec_48_T_3[5:0] ? myVec_3 : _GEN_1068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1070 = 6'h4 == _myNewVec_48_T_3[5:0] ? myVec_4 : _GEN_1069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1071 = 6'h5 == _myNewVec_48_T_3[5:0] ? myVec_5 : _GEN_1070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1072 = 6'h6 == _myNewVec_48_T_3[5:0] ? myVec_6 : _GEN_1071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1073 = 6'h7 == _myNewVec_48_T_3[5:0] ? myVec_7 : _GEN_1072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1074 = 6'h8 == _myNewVec_48_T_3[5:0] ? myVec_8 : _GEN_1073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1075 = 6'h9 == _myNewVec_48_T_3[5:0] ? myVec_9 : _GEN_1074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1076 = 6'ha == _myNewVec_48_T_3[5:0] ? myVec_10 : _GEN_1075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1077 = 6'hb == _myNewVec_48_T_3[5:0] ? myVec_11 : _GEN_1076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1078 = 6'hc == _myNewVec_48_T_3[5:0] ? myVec_12 : _GEN_1077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1079 = 6'hd == _myNewVec_48_T_3[5:0] ? myVec_13 : _GEN_1078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1080 = 6'he == _myNewVec_48_T_3[5:0] ? myVec_14 : _GEN_1079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1081 = 6'hf == _myNewVec_48_T_3[5:0] ? myVec_15 : _GEN_1080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1082 = 6'h10 == _myNewVec_48_T_3[5:0] ? myVec_16 : _GEN_1081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1083 = 6'h11 == _myNewVec_48_T_3[5:0] ? myVec_17 : _GEN_1082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1084 = 6'h12 == _myNewVec_48_T_3[5:0] ? myVec_18 : _GEN_1083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1085 = 6'h13 == _myNewVec_48_T_3[5:0] ? myVec_19 : _GEN_1084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1086 = 6'h14 == _myNewVec_48_T_3[5:0] ? myVec_20 : _GEN_1085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1087 = 6'h15 == _myNewVec_48_T_3[5:0] ? myVec_21 : _GEN_1086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1088 = 6'h16 == _myNewVec_48_T_3[5:0] ? myVec_22 : _GEN_1087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1089 = 6'h17 == _myNewVec_48_T_3[5:0] ? myVec_23 : _GEN_1088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1090 = 6'h18 == _myNewVec_48_T_3[5:0] ? myVec_24 : _GEN_1089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1091 = 6'h19 == _myNewVec_48_T_3[5:0] ? myVec_25 : _GEN_1090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1092 = 6'h1a == _myNewVec_48_T_3[5:0] ? myVec_26 : _GEN_1091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1093 = 6'h1b == _myNewVec_48_T_3[5:0] ? myVec_27 : _GEN_1092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1094 = 6'h1c == _myNewVec_48_T_3[5:0] ? myVec_28 : _GEN_1093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1095 = 6'h1d == _myNewVec_48_T_3[5:0] ? myVec_29 : _GEN_1094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1096 = 6'h1e == _myNewVec_48_T_3[5:0] ? myVec_30 : _GEN_1095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1097 = 6'h1f == _myNewVec_48_T_3[5:0] ? myVec_31 : _GEN_1096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1098 = 6'h20 == _myNewVec_48_T_3[5:0] ? myVec_32 : _GEN_1097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1099 = 6'h21 == _myNewVec_48_T_3[5:0] ? myVec_33 : _GEN_1098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1100 = 6'h22 == _myNewVec_48_T_3[5:0] ? myVec_34 : _GEN_1099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1101 = 6'h23 == _myNewVec_48_T_3[5:0] ? myVec_35 : _GEN_1100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1102 = 6'h24 == _myNewVec_48_T_3[5:0] ? myVec_36 : _GEN_1101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1103 = 6'h25 == _myNewVec_48_T_3[5:0] ? myVec_37 : _GEN_1102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1104 = 6'h26 == _myNewVec_48_T_3[5:0] ? myVec_38 : _GEN_1103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1105 = 6'h27 == _myNewVec_48_T_3[5:0] ? myVec_39 : _GEN_1104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1106 = 6'h28 == _myNewVec_48_T_3[5:0] ? myVec_40 : _GEN_1105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1107 = 6'h29 == _myNewVec_48_T_3[5:0] ? myVec_41 : _GEN_1106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1108 = 6'h2a == _myNewVec_48_T_3[5:0] ? myVec_42 : _GEN_1107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1109 = 6'h2b == _myNewVec_48_T_3[5:0] ? myVec_43 : _GEN_1108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1110 = 6'h2c == _myNewVec_48_T_3[5:0] ? myVec_44 : _GEN_1109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1111 = 6'h2d == _myNewVec_48_T_3[5:0] ? myVec_45 : _GEN_1110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1112 = 6'h2e == _myNewVec_48_T_3[5:0] ? myVec_46 : _GEN_1111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1113 = 6'h2f == _myNewVec_48_T_3[5:0] ? myVec_47 : _GEN_1112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1114 = 6'h30 == _myNewVec_48_T_3[5:0] ? myVec_48 : _GEN_1113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1115 = 6'h31 == _myNewVec_48_T_3[5:0] ? myVec_49 : _GEN_1114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1116 = 6'h32 == _myNewVec_48_T_3[5:0] ? myVec_50 : _GEN_1115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1117 = 6'h33 == _myNewVec_48_T_3[5:0] ? myVec_51 : _GEN_1116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1118 = 6'h34 == _myNewVec_48_T_3[5:0] ? myVec_52 : _GEN_1117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1119 = 6'h35 == _myNewVec_48_T_3[5:0] ? myVec_53 : _GEN_1118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1120 = 6'h36 == _myNewVec_48_T_3[5:0] ? myVec_54 : _GEN_1119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1121 = 6'h37 == _myNewVec_48_T_3[5:0] ? myVec_55 : _GEN_1120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1122 = 6'h38 == _myNewVec_48_T_3[5:0] ? myVec_56 : _GEN_1121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1123 = 6'h39 == _myNewVec_48_T_3[5:0] ? myVec_57 : _GEN_1122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1124 = 6'h3a == _myNewVec_48_T_3[5:0] ? myVec_58 : _GEN_1123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1125 = 6'h3b == _myNewVec_48_T_3[5:0] ? myVec_59 : _GEN_1124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1126 = 6'h3c == _myNewVec_48_T_3[5:0] ? myVec_60 : _GEN_1125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1127 = 6'h3d == _myNewVec_48_T_3[5:0] ? myVec_61 : _GEN_1126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1128 = 6'h3e == _myNewVec_48_T_3[5:0] ? myVec_62 : _GEN_1127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_48 = 6'h3f == _myNewVec_48_T_3[5:0] ? myVec_63 : _GEN_1128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_hi_lo = {myNewVec_55,myNewVec_54,myNewVec_53,myNewVec_52,myNewVec_51,myNewVec_50,myNewVec_49
    ,myNewVec_48}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_47_T_3 = _myNewVec_63_T_1 + 16'h10; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1131 = 6'h1 == _myNewVec_47_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1132 = 6'h2 == _myNewVec_47_T_3[5:0] ? myVec_2 : _GEN_1131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1133 = 6'h3 == _myNewVec_47_T_3[5:0] ? myVec_3 : _GEN_1132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1134 = 6'h4 == _myNewVec_47_T_3[5:0] ? myVec_4 : _GEN_1133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1135 = 6'h5 == _myNewVec_47_T_3[5:0] ? myVec_5 : _GEN_1134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1136 = 6'h6 == _myNewVec_47_T_3[5:0] ? myVec_6 : _GEN_1135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1137 = 6'h7 == _myNewVec_47_T_3[5:0] ? myVec_7 : _GEN_1136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1138 = 6'h8 == _myNewVec_47_T_3[5:0] ? myVec_8 : _GEN_1137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1139 = 6'h9 == _myNewVec_47_T_3[5:0] ? myVec_9 : _GEN_1138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1140 = 6'ha == _myNewVec_47_T_3[5:0] ? myVec_10 : _GEN_1139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1141 = 6'hb == _myNewVec_47_T_3[5:0] ? myVec_11 : _GEN_1140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1142 = 6'hc == _myNewVec_47_T_3[5:0] ? myVec_12 : _GEN_1141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1143 = 6'hd == _myNewVec_47_T_3[5:0] ? myVec_13 : _GEN_1142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1144 = 6'he == _myNewVec_47_T_3[5:0] ? myVec_14 : _GEN_1143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1145 = 6'hf == _myNewVec_47_T_3[5:0] ? myVec_15 : _GEN_1144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1146 = 6'h10 == _myNewVec_47_T_3[5:0] ? myVec_16 : _GEN_1145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1147 = 6'h11 == _myNewVec_47_T_3[5:0] ? myVec_17 : _GEN_1146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1148 = 6'h12 == _myNewVec_47_T_3[5:0] ? myVec_18 : _GEN_1147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1149 = 6'h13 == _myNewVec_47_T_3[5:0] ? myVec_19 : _GEN_1148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1150 = 6'h14 == _myNewVec_47_T_3[5:0] ? myVec_20 : _GEN_1149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1151 = 6'h15 == _myNewVec_47_T_3[5:0] ? myVec_21 : _GEN_1150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1152 = 6'h16 == _myNewVec_47_T_3[5:0] ? myVec_22 : _GEN_1151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1153 = 6'h17 == _myNewVec_47_T_3[5:0] ? myVec_23 : _GEN_1152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1154 = 6'h18 == _myNewVec_47_T_3[5:0] ? myVec_24 : _GEN_1153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1155 = 6'h19 == _myNewVec_47_T_3[5:0] ? myVec_25 : _GEN_1154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1156 = 6'h1a == _myNewVec_47_T_3[5:0] ? myVec_26 : _GEN_1155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1157 = 6'h1b == _myNewVec_47_T_3[5:0] ? myVec_27 : _GEN_1156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1158 = 6'h1c == _myNewVec_47_T_3[5:0] ? myVec_28 : _GEN_1157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1159 = 6'h1d == _myNewVec_47_T_3[5:0] ? myVec_29 : _GEN_1158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1160 = 6'h1e == _myNewVec_47_T_3[5:0] ? myVec_30 : _GEN_1159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1161 = 6'h1f == _myNewVec_47_T_3[5:0] ? myVec_31 : _GEN_1160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1162 = 6'h20 == _myNewVec_47_T_3[5:0] ? myVec_32 : _GEN_1161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1163 = 6'h21 == _myNewVec_47_T_3[5:0] ? myVec_33 : _GEN_1162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1164 = 6'h22 == _myNewVec_47_T_3[5:0] ? myVec_34 : _GEN_1163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1165 = 6'h23 == _myNewVec_47_T_3[5:0] ? myVec_35 : _GEN_1164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1166 = 6'h24 == _myNewVec_47_T_3[5:0] ? myVec_36 : _GEN_1165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1167 = 6'h25 == _myNewVec_47_T_3[5:0] ? myVec_37 : _GEN_1166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1168 = 6'h26 == _myNewVec_47_T_3[5:0] ? myVec_38 : _GEN_1167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1169 = 6'h27 == _myNewVec_47_T_3[5:0] ? myVec_39 : _GEN_1168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1170 = 6'h28 == _myNewVec_47_T_3[5:0] ? myVec_40 : _GEN_1169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1171 = 6'h29 == _myNewVec_47_T_3[5:0] ? myVec_41 : _GEN_1170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1172 = 6'h2a == _myNewVec_47_T_3[5:0] ? myVec_42 : _GEN_1171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1173 = 6'h2b == _myNewVec_47_T_3[5:0] ? myVec_43 : _GEN_1172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1174 = 6'h2c == _myNewVec_47_T_3[5:0] ? myVec_44 : _GEN_1173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1175 = 6'h2d == _myNewVec_47_T_3[5:0] ? myVec_45 : _GEN_1174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1176 = 6'h2e == _myNewVec_47_T_3[5:0] ? myVec_46 : _GEN_1175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1177 = 6'h2f == _myNewVec_47_T_3[5:0] ? myVec_47 : _GEN_1176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1178 = 6'h30 == _myNewVec_47_T_3[5:0] ? myVec_48 : _GEN_1177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1179 = 6'h31 == _myNewVec_47_T_3[5:0] ? myVec_49 : _GEN_1178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1180 = 6'h32 == _myNewVec_47_T_3[5:0] ? myVec_50 : _GEN_1179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1181 = 6'h33 == _myNewVec_47_T_3[5:0] ? myVec_51 : _GEN_1180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1182 = 6'h34 == _myNewVec_47_T_3[5:0] ? myVec_52 : _GEN_1181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1183 = 6'h35 == _myNewVec_47_T_3[5:0] ? myVec_53 : _GEN_1182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1184 = 6'h36 == _myNewVec_47_T_3[5:0] ? myVec_54 : _GEN_1183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1185 = 6'h37 == _myNewVec_47_T_3[5:0] ? myVec_55 : _GEN_1184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1186 = 6'h38 == _myNewVec_47_T_3[5:0] ? myVec_56 : _GEN_1185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1187 = 6'h39 == _myNewVec_47_T_3[5:0] ? myVec_57 : _GEN_1186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1188 = 6'h3a == _myNewVec_47_T_3[5:0] ? myVec_58 : _GEN_1187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1189 = 6'h3b == _myNewVec_47_T_3[5:0] ? myVec_59 : _GEN_1188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1190 = 6'h3c == _myNewVec_47_T_3[5:0] ? myVec_60 : _GEN_1189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1191 = 6'h3d == _myNewVec_47_T_3[5:0] ? myVec_61 : _GEN_1190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1192 = 6'h3e == _myNewVec_47_T_3[5:0] ? myVec_62 : _GEN_1191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_47 = 6'h3f == _myNewVec_47_T_3[5:0] ? myVec_63 : _GEN_1192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_46_T_3 = _myNewVec_63_T_1 + 16'h11; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1195 = 6'h1 == _myNewVec_46_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1196 = 6'h2 == _myNewVec_46_T_3[5:0] ? myVec_2 : _GEN_1195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1197 = 6'h3 == _myNewVec_46_T_3[5:0] ? myVec_3 : _GEN_1196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1198 = 6'h4 == _myNewVec_46_T_3[5:0] ? myVec_4 : _GEN_1197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1199 = 6'h5 == _myNewVec_46_T_3[5:0] ? myVec_5 : _GEN_1198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1200 = 6'h6 == _myNewVec_46_T_3[5:0] ? myVec_6 : _GEN_1199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1201 = 6'h7 == _myNewVec_46_T_3[5:0] ? myVec_7 : _GEN_1200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1202 = 6'h8 == _myNewVec_46_T_3[5:0] ? myVec_8 : _GEN_1201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1203 = 6'h9 == _myNewVec_46_T_3[5:0] ? myVec_9 : _GEN_1202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1204 = 6'ha == _myNewVec_46_T_3[5:0] ? myVec_10 : _GEN_1203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1205 = 6'hb == _myNewVec_46_T_3[5:0] ? myVec_11 : _GEN_1204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1206 = 6'hc == _myNewVec_46_T_3[5:0] ? myVec_12 : _GEN_1205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1207 = 6'hd == _myNewVec_46_T_3[5:0] ? myVec_13 : _GEN_1206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1208 = 6'he == _myNewVec_46_T_3[5:0] ? myVec_14 : _GEN_1207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1209 = 6'hf == _myNewVec_46_T_3[5:0] ? myVec_15 : _GEN_1208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1210 = 6'h10 == _myNewVec_46_T_3[5:0] ? myVec_16 : _GEN_1209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1211 = 6'h11 == _myNewVec_46_T_3[5:0] ? myVec_17 : _GEN_1210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1212 = 6'h12 == _myNewVec_46_T_3[5:0] ? myVec_18 : _GEN_1211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1213 = 6'h13 == _myNewVec_46_T_3[5:0] ? myVec_19 : _GEN_1212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1214 = 6'h14 == _myNewVec_46_T_3[5:0] ? myVec_20 : _GEN_1213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1215 = 6'h15 == _myNewVec_46_T_3[5:0] ? myVec_21 : _GEN_1214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1216 = 6'h16 == _myNewVec_46_T_3[5:0] ? myVec_22 : _GEN_1215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1217 = 6'h17 == _myNewVec_46_T_3[5:0] ? myVec_23 : _GEN_1216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1218 = 6'h18 == _myNewVec_46_T_3[5:0] ? myVec_24 : _GEN_1217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1219 = 6'h19 == _myNewVec_46_T_3[5:0] ? myVec_25 : _GEN_1218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1220 = 6'h1a == _myNewVec_46_T_3[5:0] ? myVec_26 : _GEN_1219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1221 = 6'h1b == _myNewVec_46_T_3[5:0] ? myVec_27 : _GEN_1220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1222 = 6'h1c == _myNewVec_46_T_3[5:0] ? myVec_28 : _GEN_1221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1223 = 6'h1d == _myNewVec_46_T_3[5:0] ? myVec_29 : _GEN_1222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1224 = 6'h1e == _myNewVec_46_T_3[5:0] ? myVec_30 : _GEN_1223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1225 = 6'h1f == _myNewVec_46_T_3[5:0] ? myVec_31 : _GEN_1224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1226 = 6'h20 == _myNewVec_46_T_3[5:0] ? myVec_32 : _GEN_1225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1227 = 6'h21 == _myNewVec_46_T_3[5:0] ? myVec_33 : _GEN_1226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1228 = 6'h22 == _myNewVec_46_T_3[5:0] ? myVec_34 : _GEN_1227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1229 = 6'h23 == _myNewVec_46_T_3[5:0] ? myVec_35 : _GEN_1228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1230 = 6'h24 == _myNewVec_46_T_3[5:0] ? myVec_36 : _GEN_1229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1231 = 6'h25 == _myNewVec_46_T_3[5:0] ? myVec_37 : _GEN_1230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1232 = 6'h26 == _myNewVec_46_T_3[5:0] ? myVec_38 : _GEN_1231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1233 = 6'h27 == _myNewVec_46_T_3[5:0] ? myVec_39 : _GEN_1232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1234 = 6'h28 == _myNewVec_46_T_3[5:0] ? myVec_40 : _GEN_1233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1235 = 6'h29 == _myNewVec_46_T_3[5:0] ? myVec_41 : _GEN_1234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1236 = 6'h2a == _myNewVec_46_T_3[5:0] ? myVec_42 : _GEN_1235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1237 = 6'h2b == _myNewVec_46_T_3[5:0] ? myVec_43 : _GEN_1236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1238 = 6'h2c == _myNewVec_46_T_3[5:0] ? myVec_44 : _GEN_1237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1239 = 6'h2d == _myNewVec_46_T_3[5:0] ? myVec_45 : _GEN_1238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1240 = 6'h2e == _myNewVec_46_T_3[5:0] ? myVec_46 : _GEN_1239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1241 = 6'h2f == _myNewVec_46_T_3[5:0] ? myVec_47 : _GEN_1240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1242 = 6'h30 == _myNewVec_46_T_3[5:0] ? myVec_48 : _GEN_1241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1243 = 6'h31 == _myNewVec_46_T_3[5:0] ? myVec_49 : _GEN_1242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1244 = 6'h32 == _myNewVec_46_T_3[5:0] ? myVec_50 : _GEN_1243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1245 = 6'h33 == _myNewVec_46_T_3[5:0] ? myVec_51 : _GEN_1244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1246 = 6'h34 == _myNewVec_46_T_3[5:0] ? myVec_52 : _GEN_1245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1247 = 6'h35 == _myNewVec_46_T_3[5:0] ? myVec_53 : _GEN_1246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1248 = 6'h36 == _myNewVec_46_T_3[5:0] ? myVec_54 : _GEN_1247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1249 = 6'h37 == _myNewVec_46_T_3[5:0] ? myVec_55 : _GEN_1248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1250 = 6'h38 == _myNewVec_46_T_3[5:0] ? myVec_56 : _GEN_1249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1251 = 6'h39 == _myNewVec_46_T_3[5:0] ? myVec_57 : _GEN_1250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1252 = 6'h3a == _myNewVec_46_T_3[5:0] ? myVec_58 : _GEN_1251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1253 = 6'h3b == _myNewVec_46_T_3[5:0] ? myVec_59 : _GEN_1252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1254 = 6'h3c == _myNewVec_46_T_3[5:0] ? myVec_60 : _GEN_1253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1255 = 6'h3d == _myNewVec_46_T_3[5:0] ? myVec_61 : _GEN_1254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1256 = 6'h3e == _myNewVec_46_T_3[5:0] ? myVec_62 : _GEN_1255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_46 = 6'h3f == _myNewVec_46_T_3[5:0] ? myVec_63 : _GEN_1256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_45_T_3 = _myNewVec_63_T_1 + 16'h12; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1259 = 6'h1 == _myNewVec_45_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1260 = 6'h2 == _myNewVec_45_T_3[5:0] ? myVec_2 : _GEN_1259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1261 = 6'h3 == _myNewVec_45_T_3[5:0] ? myVec_3 : _GEN_1260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1262 = 6'h4 == _myNewVec_45_T_3[5:0] ? myVec_4 : _GEN_1261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1263 = 6'h5 == _myNewVec_45_T_3[5:0] ? myVec_5 : _GEN_1262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1264 = 6'h6 == _myNewVec_45_T_3[5:0] ? myVec_6 : _GEN_1263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1265 = 6'h7 == _myNewVec_45_T_3[5:0] ? myVec_7 : _GEN_1264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1266 = 6'h8 == _myNewVec_45_T_3[5:0] ? myVec_8 : _GEN_1265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1267 = 6'h9 == _myNewVec_45_T_3[5:0] ? myVec_9 : _GEN_1266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1268 = 6'ha == _myNewVec_45_T_3[5:0] ? myVec_10 : _GEN_1267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1269 = 6'hb == _myNewVec_45_T_3[5:0] ? myVec_11 : _GEN_1268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1270 = 6'hc == _myNewVec_45_T_3[5:0] ? myVec_12 : _GEN_1269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1271 = 6'hd == _myNewVec_45_T_3[5:0] ? myVec_13 : _GEN_1270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1272 = 6'he == _myNewVec_45_T_3[5:0] ? myVec_14 : _GEN_1271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1273 = 6'hf == _myNewVec_45_T_3[5:0] ? myVec_15 : _GEN_1272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1274 = 6'h10 == _myNewVec_45_T_3[5:0] ? myVec_16 : _GEN_1273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1275 = 6'h11 == _myNewVec_45_T_3[5:0] ? myVec_17 : _GEN_1274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1276 = 6'h12 == _myNewVec_45_T_3[5:0] ? myVec_18 : _GEN_1275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1277 = 6'h13 == _myNewVec_45_T_3[5:0] ? myVec_19 : _GEN_1276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1278 = 6'h14 == _myNewVec_45_T_3[5:0] ? myVec_20 : _GEN_1277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1279 = 6'h15 == _myNewVec_45_T_3[5:0] ? myVec_21 : _GEN_1278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1280 = 6'h16 == _myNewVec_45_T_3[5:0] ? myVec_22 : _GEN_1279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1281 = 6'h17 == _myNewVec_45_T_3[5:0] ? myVec_23 : _GEN_1280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1282 = 6'h18 == _myNewVec_45_T_3[5:0] ? myVec_24 : _GEN_1281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1283 = 6'h19 == _myNewVec_45_T_3[5:0] ? myVec_25 : _GEN_1282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1284 = 6'h1a == _myNewVec_45_T_3[5:0] ? myVec_26 : _GEN_1283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1285 = 6'h1b == _myNewVec_45_T_3[5:0] ? myVec_27 : _GEN_1284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1286 = 6'h1c == _myNewVec_45_T_3[5:0] ? myVec_28 : _GEN_1285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1287 = 6'h1d == _myNewVec_45_T_3[5:0] ? myVec_29 : _GEN_1286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1288 = 6'h1e == _myNewVec_45_T_3[5:0] ? myVec_30 : _GEN_1287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1289 = 6'h1f == _myNewVec_45_T_3[5:0] ? myVec_31 : _GEN_1288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1290 = 6'h20 == _myNewVec_45_T_3[5:0] ? myVec_32 : _GEN_1289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1291 = 6'h21 == _myNewVec_45_T_3[5:0] ? myVec_33 : _GEN_1290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1292 = 6'h22 == _myNewVec_45_T_3[5:0] ? myVec_34 : _GEN_1291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1293 = 6'h23 == _myNewVec_45_T_3[5:0] ? myVec_35 : _GEN_1292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1294 = 6'h24 == _myNewVec_45_T_3[5:0] ? myVec_36 : _GEN_1293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1295 = 6'h25 == _myNewVec_45_T_3[5:0] ? myVec_37 : _GEN_1294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1296 = 6'h26 == _myNewVec_45_T_3[5:0] ? myVec_38 : _GEN_1295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1297 = 6'h27 == _myNewVec_45_T_3[5:0] ? myVec_39 : _GEN_1296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1298 = 6'h28 == _myNewVec_45_T_3[5:0] ? myVec_40 : _GEN_1297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1299 = 6'h29 == _myNewVec_45_T_3[5:0] ? myVec_41 : _GEN_1298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1300 = 6'h2a == _myNewVec_45_T_3[5:0] ? myVec_42 : _GEN_1299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1301 = 6'h2b == _myNewVec_45_T_3[5:0] ? myVec_43 : _GEN_1300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1302 = 6'h2c == _myNewVec_45_T_3[5:0] ? myVec_44 : _GEN_1301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1303 = 6'h2d == _myNewVec_45_T_3[5:0] ? myVec_45 : _GEN_1302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1304 = 6'h2e == _myNewVec_45_T_3[5:0] ? myVec_46 : _GEN_1303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1305 = 6'h2f == _myNewVec_45_T_3[5:0] ? myVec_47 : _GEN_1304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1306 = 6'h30 == _myNewVec_45_T_3[5:0] ? myVec_48 : _GEN_1305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1307 = 6'h31 == _myNewVec_45_T_3[5:0] ? myVec_49 : _GEN_1306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1308 = 6'h32 == _myNewVec_45_T_3[5:0] ? myVec_50 : _GEN_1307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1309 = 6'h33 == _myNewVec_45_T_3[5:0] ? myVec_51 : _GEN_1308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1310 = 6'h34 == _myNewVec_45_T_3[5:0] ? myVec_52 : _GEN_1309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1311 = 6'h35 == _myNewVec_45_T_3[5:0] ? myVec_53 : _GEN_1310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1312 = 6'h36 == _myNewVec_45_T_3[5:0] ? myVec_54 : _GEN_1311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1313 = 6'h37 == _myNewVec_45_T_3[5:0] ? myVec_55 : _GEN_1312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1314 = 6'h38 == _myNewVec_45_T_3[5:0] ? myVec_56 : _GEN_1313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1315 = 6'h39 == _myNewVec_45_T_3[5:0] ? myVec_57 : _GEN_1314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1316 = 6'h3a == _myNewVec_45_T_3[5:0] ? myVec_58 : _GEN_1315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1317 = 6'h3b == _myNewVec_45_T_3[5:0] ? myVec_59 : _GEN_1316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1318 = 6'h3c == _myNewVec_45_T_3[5:0] ? myVec_60 : _GEN_1317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1319 = 6'h3d == _myNewVec_45_T_3[5:0] ? myVec_61 : _GEN_1318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1320 = 6'h3e == _myNewVec_45_T_3[5:0] ? myVec_62 : _GEN_1319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_45 = 6'h3f == _myNewVec_45_T_3[5:0] ? myVec_63 : _GEN_1320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_44_T_3 = _myNewVec_63_T_1 + 16'h13; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1323 = 6'h1 == _myNewVec_44_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1324 = 6'h2 == _myNewVec_44_T_3[5:0] ? myVec_2 : _GEN_1323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1325 = 6'h3 == _myNewVec_44_T_3[5:0] ? myVec_3 : _GEN_1324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1326 = 6'h4 == _myNewVec_44_T_3[5:0] ? myVec_4 : _GEN_1325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1327 = 6'h5 == _myNewVec_44_T_3[5:0] ? myVec_5 : _GEN_1326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1328 = 6'h6 == _myNewVec_44_T_3[5:0] ? myVec_6 : _GEN_1327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1329 = 6'h7 == _myNewVec_44_T_3[5:0] ? myVec_7 : _GEN_1328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1330 = 6'h8 == _myNewVec_44_T_3[5:0] ? myVec_8 : _GEN_1329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1331 = 6'h9 == _myNewVec_44_T_3[5:0] ? myVec_9 : _GEN_1330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1332 = 6'ha == _myNewVec_44_T_3[5:0] ? myVec_10 : _GEN_1331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1333 = 6'hb == _myNewVec_44_T_3[5:0] ? myVec_11 : _GEN_1332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1334 = 6'hc == _myNewVec_44_T_3[5:0] ? myVec_12 : _GEN_1333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1335 = 6'hd == _myNewVec_44_T_3[5:0] ? myVec_13 : _GEN_1334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1336 = 6'he == _myNewVec_44_T_3[5:0] ? myVec_14 : _GEN_1335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1337 = 6'hf == _myNewVec_44_T_3[5:0] ? myVec_15 : _GEN_1336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1338 = 6'h10 == _myNewVec_44_T_3[5:0] ? myVec_16 : _GEN_1337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1339 = 6'h11 == _myNewVec_44_T_3[5:0] ? myVec_17 : _GEN_1338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1340 = 6'h12 == _myNewVec_44_T_3[5:0] ? myVec_18 : _GEN_1339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1341 = 6'h13 == _myNewVec_44_T_3[5:0] ? myVec_19 : _GEN_1340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1342 = 6'h14 == _myNewVec_44_T_3[5:0] ? myVec_20 : _GEN_1341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1343 = 6'h15 == _myNewVec_44_T_3[5:0] ? myVec_21 : _GEN_1342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1344 = 6'h16 == _myNewVec_44_T_3[5:0] ? myVec_22 : _GEN_1343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1345 = 6'h17 == _myNewVec_44_T_3[5:0] ? myVec_23 : _GEN_1344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1346 = 6'h18 == _myNewVec_44_T_3[5:0] ? myVec_24 : _GEN_1345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1347 = 6'h19 == _myNewVec_44_T_3[5:0] ? myVec_25 : _GEN_1346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1348 = 6'h1a == _myNewVec_44_T_3[5:0] ? myVec_26 : _GEN_1347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1349 = 6'h1b == _myNewVec_44_T_3[5:0] ? myVec_27 : _GEN_1348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1350 = 6'h1c == _myNewVec_44_T_3[5:0] ? myVec_28 : _GEN_1349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1351 = 6'h1d == _myNewVec_44_T_3[5:0] ? myVec_29 : _GEN_1350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1352 = 6'h1e == _myNewVec_44_T_3[5:0] ? myVec_30 : _GEN_1351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1353 = 6'h1f == _myNewVec_44_T_3[5:0] ? myVec_31 : _GEN_1352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1354 = 6'h20 == _myNewVec_44_T_3[5:0] ? myVec_32 : _GEN_1353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1355 = 6'h21 == _myNewVec_44_T_3[5:0] ? myVec_33 : _GEN_1354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1356 = 6'h22 == _myNewVec_44_T_3[5:0] ? myVec_34 : _GEN_1355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1357 = 6'h23 == _myNewVec_44_T_3[5:0] ? myVec_35 : _GEN_1356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1358 = 6'h24 == _myNewVec_44_T_3[5:0] ? myVec_36 : _GEN_1357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1359 = 6'h25 == _myNewVec_44_T_3[5:0] ? myVec_37 : _GEN_1358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1360 = 6'h26 == _myNewVec_44_T_3[5:0] ? myVec_38 : _GEN_1359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1361 = 6'h27 == _myNewVec_44_T_3[5:0] ? myVec_39 : _GEN_1360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1362 = 6'h28 == _myNewVec_44_T_3[5:0] ? myVec_40 : _GEN_1361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1363 = 6'h29 == _myNewVec_44_T_3[5:0] ? myVec_41 : _GEN_1362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1364 = 6'h2a == _myNewVec_44_T_3[5:0] ? myVec_42 : _GEN_1363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1365 = 6'h2b == _myNewVec_44_T_3[5:0] ? myVec_43 : _GEN_1364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1366 = 6'h2c == _myNewVec_44_T_3[5:0] ? myVec_44 : _GEN_1365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1367 = 6'h2d == _myNewVec_44_T_3[5:0] ? myVec_45 : _GEN_1366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1368 = 6'h2e == _myNewVec_44_T_3[5:0] ? myVec_46 : _GEN_1367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1369 = 6'h2f == _myNewVec_44_T_3[5:0] ? myVec_47 : _GEN_1368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1370 = 6'h30 == _myNewVec_44_T_3[5:0] ? myVec_48 : _GEN_1369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1371 = 6'h31 == _myNewVec_44_T_3[5:0] ? myVec_49 : _GEN_1370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1372 = 6'h32 == _myNewVec_44_T_3[5:0] ? myVec_50 : _GEN_1371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1373 = 6'h33 == _myNewVec_44_T_3[5:0] ? myVec_51 : _GEN_1372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1374 = 6'h34 == _myNewVec_44_T_3[5:0] ? myVec_52 : _GEN_1373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1375 = 6'h35 == _myNewVec_44_T_3[5:0] ? myVec_53 : _GEN_1374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1376 = 6'h36 == _myNewVec_44_T_3[5:0] ? myVec_54 : _GEN_1375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1377 = 6'h37 == _myNewVec_44_T_3[5:0] ? myVec_55 : _GEN_1376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1378 = 6'h38 == _myNewVec_44_T_3[5:0] ? myVec_56 : _GEN_1377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1379 = 6'h39 == _myNewVec_44_T_3[5:0] ? myVec_57 : _GEN_1378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1380 = 6'h3a == _myNewVec_44_T_3[5:0] ? myVec_58 : _GEN_1379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1381 = 6'h3b == _myNewVec_44_T_3[5:0] ? myVec_59 : _GEN_1380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1382 = 6'h3c == _myNewVec_44_T_3[5:0] ? myVec_60 : _GEN_1381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1383 = 6'h3d == _myNewVec_44_T_3[5:0] ? myVec_61 : _GEN_1382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1384 = 6'h3e == _myNewVec_44_T_3[5:0] ? myVec_62 : _GEN_1383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_44 = 6'h3f == _myNewVec_44_T_3[5:0] ? myVec_63 : _GEN_1384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_43_T_3 = _myNewVec_63_T_1 + 16'h14; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1387 = 6'h1 == _myNewVec_43_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1388 = 6'h2 == _myNewVec_43_T_3[5:0] ? myVec_2 : _GEN_1387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1389 = 6'h3 == _myNewVec_43_T_3[5:0] ? myVec_3 : _GEN_1388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1390 = 6'h4 == _myNewVec_43_T_3[5:0] ? myVec_4 : _GEN_1389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1391 = 6'h5 == _myNewVec_43_T_3[5:0] ? myVec_5 : _GEN_1390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1392 = 6'h6 == _myNewVec_43_T_3[5:0] ? myVec_6 : _GEN_1391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1393 = 6'h7 == _myNewVec_43_T_3[5:0] ? myVec_7 : _GEN_1392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1394 = 6'h8 == _myNewVec_43_T_3[5:0] ? myVec_8 : _GEN_1393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1395 = 6'h9 == _myNewVec_43_T_3[5:0] ? myVec_9 : _GEN_1394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1396 = 6'ha == _myNewVec_43_T_3[5:0] ? myVec_10 : _GEN_1395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1397 = 6'hb == _myNewVec_43_T_3[5:0] ? myVec_11 : _GEN_1396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1398 = 6'hc == _myNewVec_43_T_3[5:0] ? myVec_12 : _GEN_1397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1399 = 6'hd == _myNewVec_43_T_3[5:0] ? myVec_13 : _GEN_1398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1400 = 6'he == _myNewVec_43_T_3[5:0] ? myVec_14 : _GEN_1399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1401 = 6'hf == _myNewVec_43_T_3[5:0] ? myVec_15 : _GEN_1400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1402 = 6'h10 == _myNewVec_43_T_3[5:0] ? myVec_16 : _GEN_1401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1403 = 6'h11 == _myNewVec_43_T_3[5:0] ? myVec_17 : _GEN_1402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1404 = 6'h12 == _myNewVec_43_T_3[5:0] ? myVec_18 : _GEN_1403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1405 = 6'h13 == _myNewVec_43_T_3[5:0] ? myVec_19 : _GEN_1404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1406 = 6'h14 == _myNewVec_43_T_3[5:0] ? myVec_20 : _GEN_1405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1407 = 6'h15 == _myNewVec_43_T_3[5:0] ? myVec_21 : _GEN_1406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1408 = 6'h16 == _myNewVec_43_T_3[5:0] ? myVec_22 : _GEN_1407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1409 = 6'h17 == _myNewVec_43_T_3[5:0] ? myVec_23 : _GEN_1408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1410 = 6'h18 == _myNewVec_43_T_3[5:0] ? myVec_24 : _GEN_1409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1411 = 6'h19 == _myNewVec_43_T_3[5:0] ? myVec_25 : _GEN_1410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1412 = 6'h1a == _myNewVec_43_T_3[5:0] ? myVec_26 : _GEN_1411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1413 = 6'h1b == _myNewVec_43_T_3[5:0] ? myVec_27 : _GEN_1412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1414 = 6'h1c == _myNewVec_43_T_3[5:0] ? myVec_28 : _GEN_1413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1415 = 6'h1d == _myNewVec_43_T_3[5:0] ? myVec_29 : _GEN_1414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1416 = 6'h1e == _myNewVec_43_T_3[5:0] ? myVec_30 : _GEN_1415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1417 = 6'h1f == _myNewVec_43_T_3[5:0] ? myVec_31 : _GEN_1416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1418 = 6'h20 == _myNewVec_43_T_3[5:0] ? myVec_32 : _GEN_1417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1419 = 6'h21 == _myNewVec_43_T_3[5:0] ? myVec_33 : _GEN_1418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1420 = 6'h22 == _myNewVec_43_T_3[5:0] ? myVec_34 : _GEN_1419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1421 = 6'h23 == _myNewVec_43_T_3[5:0] ? myVec_35 : _GEN_1420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1422 = 6'h24 == _myNewVec_43_T_3[5:0] ? myVec_36 : _GEN_1421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1423 = 6'h25 == _myNewVec_43_T_3[5:0] ? myVec_37 : _GEN_1422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1424 = 6'h26 == _myNewVec_43_T_3[5:0] ? myVec_38 : _GEN_1423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1425 = 6'h27 == _myNewVec_43_T_3[5:0] ? myVec_39 : _GEN_1424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1426 = 6'h28 == _myNewVec_43_T_3[5:0] ? myVec_40 : _GEN_1425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1427 = 6'h29 == _myNewVec_43_T_3[5:0] ? myVec_41 : _GEN_1426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1428 = 6'h2a == _myNewVec_43_T_3[5:0] ? myVec_42 : _GEN_1427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1429 = 6'h2b == _myNewVec_43_T_3[5:0] ? myVec_43 : _GEN_1428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1430 = 6'h2c == _myNewVec_43_T_3[5:0] ? myVec_44 : _GEN_1429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1431 = 6'h2d == _myNewVec_43_T_3[5:0] ? myVec_45 : _GEN_1430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1432 = 6'h2e == _myNewVec_43_T_3[5:0] ? myVec_46 : _GEN_1431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1433 = 6'h2f == _myNewVec_43_T_3[5:0] ? myVec_47 : _GEN_1432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1434 = 6'h30 == _myNewVec_43_T_3[5:0] ? myVec_48 : _GEN_1433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1435 = 6'h31 == _myNewVec_43_T_3[5:0] ? myVec_49 : _GEN_1434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1436 = 6'h32 == _myNewVec_43_T_3[5:0] ? myVec_50 : _GEN_1435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1437 = 6'h33 == _myNewVec_43_T_3[5:0] ? myVec_51 : _GEN_1436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1438 = 6'h34 == _myNewVec_43_T_3[5:0] ? myVec_52 : _GEN_1437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1439 = 6'h35 == _myNewVec_43_T_3[5:0] ? myVec_53 : _GEN_1438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1440 = 6'h36 == _myNewVec_43_T_3[5:0] ? myVec_54 : _GEN_1439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1441 = 6'h37 == _myNewVec_43_T_3[5:0] ? myVec_55 : _GEN_1440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1442 = 6'h38 == _myNewVec_43_T_3[5:0] ? myVec_56 : _GEN_1441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1443 = 6'h39 == _myNewVec_43_T_3[5:0] ? myVec_57 : _GEN_1442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1444 = 6'h3a == _myNewVec_43_T_3[5:0] ? myVec_58 : _GEN_1443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1445 = 6'h3b == _myNewVec_43_T_3[5:0] ? myVec_59 : _GEN_1444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1446 = 6'h3c == _myNewVec_43_T_3[5:0] ? myVec_60 : _GEN_1445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1447 = 6'h3d == _myNewVec_43_T_3[5:0] ? myVec_61 : _GEN_1446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1448 = 6'h3e == _myNewVec_43_T_3[5:0] ? myVec_62 : _GEN_1447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_43 = 6'h3f == _myNewVec_43_T_3[5:0] ? myVec_63 : _GEN_1448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_42_T_3 = _myNewVec_63_T_1 + 16'h15; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1451 = 6'h1 == _myNewVec_42_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1452 = 6'h2 == _myNewVec_42_T_3[5:0] ? myVec_2 : _GEN_1451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1453 = 6'h3 == _myNewVec_42_T_3[5:0] ? myVec_3 : _GEN_1452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1454 = 6'h4 == _myNewVec_42_T_3[5:0] ? myVec_4 : _GEN_1453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1455 = 6'h5 == _myNewVec_42_T_3[5:0] ? myVec_5 : _GEN_1454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1456 = 6'h6 == _myNewVec_42_T_3[5:0] ? myVec_6 : _GEN_1455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1457 = 6'h7 == _myNewVec_42_T_3[5:0] ? myVec_7 : _GEN_1456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1458 = 6'h8 == _myNewVec_42_T_3[5:0] ? myVec_8 : _GEN_1457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1459 = 6'h9 == _myNewVec_42_T_3[5:0] ? myVec_9 : _GEN_1458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1460 = 6'ha == _myNewVec_42_T_3[5:0] ? myVec_10 : _GEN_1459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1461 = 6'hb == _myNewVec_42_T_3[5:0] ? myVec_11 : _GEN_1460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1462 = 6'hc == _myNewVec_42_T_3[5:0] ? myVec_12 : _GEN_1461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1463 = 6'hd == _myNewVec_42_T_3[5:0] ? myVec_13 : _GEN_1462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1464 = 6'he == _myNewVec_42_T_3[5:0] ? myVec_14 : _GEN_1463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1465 = 6'hf == _myNewVec_42_T_3[5:0] ? myVec_15 : _GEN_1464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1466 = 6'h10 == _myNewVec_42_T_3[5:0] ? myVec_16 : _GEN_1465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1467 = 6'h11 == _myNewVec_42_T_3[5:0] ? myVec_17 : _GEN_1466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1468 = 6'h12 == _myNewVec_42_T_3[5:0] ? myVec_18 : _GEN_1467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1469 = 6'h13 == _myNewVec_42_T_3[5:0] ? myVec_19 : _GEN_1468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1470 = 6'h14 == _myNewVec_42_T_3[5:0] ? myVec_20 : _GEN_1469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1471 = 6'h15 == _myNewVec_42_T_3[5:0] ? myVec_21 : _GEN_1470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1472 = 6'h16 == _myNewVec_42_T_3[5:0] ? myVec_22 : _GEN_1471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1473 = 6'h17 == _myNewVec_42_T_3[5:0] ? myVec_23 : _GEN_1472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1474 = 6'h18 == _myNewVec_42_T_3[5:0] ? myVec_24 : _GEN_1473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1475 = 6'h19 == _myNewVec_42_T_3[5:0] ? myVec_25 : _GEN_1474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1476 = 6'h1a == _myNewVec_42_T_3[5:0] ? myVec_26 : _GEN_1475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1477 = 6'h1b == _myNewVec_42_T_3[5:0] ? myVec_27 : _GEN_1476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1478 = 6'h1c == _myNewVec_42_T_3[5:0] ? myVec_28 : _GEN_1477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1479 = 6'h1d == _myNewVec_42_T_3[5:0] ? myVec_29 : _GEN_1478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1480 = 6'h1e == _myNewVec_42_T_3[5:0] ? myVec_30 : _GEN_1479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1481 = 6'h1f == _myNewVec_42_T_3[5:0] ? myVec_31 : _GEN_1480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1482 = 6'h20 == _myNewVec_42_T_3[5:0] ? myVec_32 : _GEN_1481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1483 = 6'h21 == _myNewVec_42_T_3[5:0] ? myVec_33 : _GEN_1482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1484 = 6'h22 == _myNewVec_42_T_3[5:0] ? myVec_34 : _GEN_1483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1485 = 6'h23 == _myNewVec_42_T_3[5:0] ? myVec_35 : _GEN_1484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1486 = 6'h24 == _myNewVec_42_T_3[5:0] ? myVec_36 : _GEN_1485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1487 = 6'h25 == _myNewVec_42_T_3[5:0] ? myVec_37 : _GEN_1486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1488 = 6'h26 == _myNewVec_42_T_3[5:0] ? myVec_38 : _GEN_1487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1489 = 6'h27 == _myNewVec_42_T_3[5:0] ? myVec_39 : _GEN_1488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1490 = 6'h28 == _myNewVec_42_T_3[5:0] ? myVec_40 : _GEN_1489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1491 = 6'h29 == _myNewVec_42_T_3[5:0] ? myVec_41 : _GEN_1490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1492 = 6'h2a == _myNewVec_42_T_3[5:0] ? myVec_42 : _GEN_1491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1493 = 6'h2b == _myNewVec_42_T_3[5:0] ? myVec_43 : _GEN_1492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1494 = 6'h2c == _myNewVec_42_T_3[5:0] ? myVec_44 : _GEN_1493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1495 = 6'h2d == _myNewVec_42_T_3[5:0] ? myVec_45 : _GEN_1494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1496 = 6'h2e == _myNewVec_42_T_3[5:0] ? myVec_46 : _GEN_1495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1497 = 6'h2f == _myNewVec_42_T_3[5:0] ? myVec_47 : _GEN_1496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1498 = 6'h30 == _myNewVec_42_T_3[5:0] ? myVec_48 : _GEN_1497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1499 = 6'h31 == _myNewVec_42_T_3[5:0] ? myVec_49 : _GEN_1498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1500 = 6'h32 == _myNewVec_42_T_3[5:0] ? myVec_50 : _GEN_1499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1501 = 6'h33 == _myNewVec_42_T_3[5:0] ? myVec_51 : _GEN_1500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1502 = 6'h34 == _myNewVec_42_T_3[5:0] ? myVec_52 : _GEN_1501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1503 = 6'h35 == _myNewVec_42_T_3[5:0] ? myVec_53 : _GEN_1502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1504 = 6'h36 == _myNewVec_42_T_3[5:0] ? myVec_54 : _GEN_1503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1505 = 6'h37 == _myNewVec_42_T_3[5:0] ? myVec_55 : _GEN_1504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1506 = 6'h38 == _myNewVec_42_T_3[5:0] ? myVec_56 : _GEN_1505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1507 = 6'h39 == _myNewVec_42_T_3[5:0] ? myVec_57 : _GEN_1506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1508 = 6'h3a == _myNewVec_42_T_3[5:0] ? myVec_58 : _GEN_1507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1509 = 6'h3b == _myNewVec_42_T_3[5:0] ? myVec_59 : _GEN_1508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1510 = 6'h3c == _myNewVec_42_T_3[5:0] ? myVec_60 : _GEN_1509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1511 = 6'h3d == _myNewVec_42_T_3[5:0] ? myVec_61 : _GEN_1510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1512 = 6'h3e == _myNewVec_42_T_3[5:0] ? myVec_62 : _GEN_1511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_42 = 6'h3f == _myNewVec_42_T_3[5:0] ? myVec_63 : _GEN_1512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_41_T_3 = _myNewVec_63_T_1 + 16'h16; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1515 = 6'h1 == _myNewVec_41_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1516 = 6'h2 == _myNewVec_41_T_3[5:0] ? myVec_2 : _GEN_1515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1517 = 6'h3 == _myNewVec_41_T_3[5:0] ? myVec_3 : _GEN_1516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1518 = 6'h4 == _myNewVec_41_T_3[5:0] ? myVec_4 : _GEN_1517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1519 = 6'h5 == _myNewVec_41_T_3[5:0] ? myVec_5 : _GEN_1518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1520 = 6'h6 == _myNewVec_41_T_3[5:0] ? myVec_6 : _GEN_1519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1521 = 6'h7 == _myNewVec_41_T_3[5:0] ? myVec_7 : _GEN_1520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1522 = 6'h8 == _myNewVec_41_T_3[5:0] ? myVec_8 : _GEN_1521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1523 = 6'h9 == _myNewVec_41_T_3[5:0] ? myVec_9 : _GEN_1522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1524 = 6'ha == _myNewVec_41_T_3[5:0] ? myVec_10 : _GEN_1523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1525 = 6'hb == _myNewVec_41_T_3[5:0] ? myVec_11 : _GEN_1524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1526 = 6'hc == _myNewVec_41_T_3[5:0] ? myVec_12 : _GEN_1525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1527 = 6'hd == _myNewVec_41_T_3[5:0] ? myVec_13 : _GEN_1526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1528 = 6'he == _myNewVec_41_T_3[5:0] ? myVec_14 : _GEN_1527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1529 = 6'hf == _myNewVec_41_T_3[5:0] ? myVec_15 : _GEN_1528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1530 = 6'h10 == _myNewVec_41_T_3[5:0] ? myVec_16 : _GEN_1529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1531 = 6'h11 == _myNewVec_41_T_3[5:0] ? myVec_17 : _GEN_1530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1532 = 6'h12 == _myNewVec_41_T_3[5:0] ? myVec_18 : _GEN_1531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1533 = 6'h13 == _myNewVec_41_T_3[5:0] ? myVec_19 : _GEN_1532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1534 = 6'h14 == _myNewVec_41_T_3[5:0] ? myVec_20 : _GEN_1533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1535 = 6'h15 == _myNewVec_41_T_3[5:0] ? myVec_21 : _GEN_1534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1536 = 6'h16 == _myNewVec_41_T_3[5:0] ? myVec_22 : _GEN_1535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1537 = 6'h17 == _myNewVec_41_T_3[5:0] ? myVec_23 : _GEN_1536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1538 = 6'h18 == _myNewVec_41_T_3[5:0] ? myVec_24 : _GEN_1537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1539 = 6'h19 == _myNewVec_41_T_3[5:0] ? myVec_25 : _GEN_1538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1540 = 6'h1a == _myNewVec_41_T_3[5:0] ? myVec_26 : _GEN_1539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1541 = 6'h1b == _myNewVec_41_T_3[5:0] ? myVec_27 : _GEN_1540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1542 = 6'h1c == _myNewVec_41_T_3[5:0] ? myVec_28 : _GEN_1541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1543 = 6'h1d == _myNewVec_41_T_3[5:0] ? myVec_29 : _GEN_1542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1544 = 6'h1e == _myNewVec_41_T_3[5:0] ? myVec_30 : _GEN_1543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1545 = 6'h1f == _myNewVec_41_T_3[5:0] ? myVec_31 : _GEN_1544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1546 = 6'h20 == _myNewVec_41_T_3[5:0] ? myVec_32 : _GEN_1545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1547 = 6'h21 == _myNewVec_41_T_3[5:0] ? myVec_33 : _GEN_1546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1548 = 6'h22 == _myNewVec_41_T_3[5:0] ? myVec_34 : _GEN_1547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1549 = 6'h23 == _myNewVec_41_T_3[5:0] ? myVec_35 : _GEN_1548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1550 = 6'h24 == _myNewVec_41_T_3[5:0] ? myVec_36 : _GEN_1549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1551 = 6'h25 == _myNewVec_41_T_3[5:0] ? myVec_37 : _GEN_1550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1552 = 6'h26 == _myNewVec_41_T_3[5:0] ? myVec_38 : _GEN_1551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1553 = 6'h27 == _myNewVec_41_T_3[5:0] ? myVec_39 : _GEN_1552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1554 = 6'h28 == _myNewVec_41_T_3[5:0] ? myVec_40 : _GEN_1553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1555 = 6'h29 == _myNewVec_41_T_3[5:0] ? myVec_41 : _GEN_1554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1556 = 6'h2a == _myNewVec_41_T_3[5:0] ? myVec_42 : _GEN_1555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1557 = 6'h2b == _myNewVec_41_T_3[5:0] ? myVec_43 : _GEN_1556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1558 = 6'h2c == _myNewVec_41_T_3[5:0] ? myVec_44 : _GEN_1557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1559 = 6'h2d == _myNewVec_41_T_3[5:0] ? myVec_45 : _GEN_1558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1560 = 6'h2e == _myNewVec_41_T_3[5:0] ? myVec_46 : _GEN_1559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1561 = 6'h2f == _myNewVec_41_T_3[5:0] ? myVec_47 : _GEN_1560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1562 = 6'h30 == _myNewVec_41_T_3[5:0] ? myVec_48 : _GEN_1561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1563 = 6'h31 == _myNewVec_41_T_3[5:0] ? myVec_49 : _GEN_1562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1564 = 6'h32 == _myNewVec_41_T_3[5:0] ? myVec_50 : _GEN_1563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1565 = 6'h33 == _myNewVec_41_T_3[5:0] ? myVec_51 : _GEN_1564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1566 = 6'h34 == _myNewVec_41_T_3[5:0] ? myVec_52 : _GEN_1565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1567 = 6'h35 == _myNewVec_41_T_3[5:0] ? myVec_53 : _GEN_1566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1568 = 6'h36 == _myNewVec_41_T_3[5:0] ? myVec_54 : _GEN_1567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1569 = 6'h37 == _myNewVec_41_T_3[5:0] ? myVec_55 : _GEN_1568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1570 = 6'h38 == _myNewVec_41_T_3[5:0] ? myVec_56 : _GEN_1569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1571 = 6'h39 == _myNewVec_41_T_3[5:0] ? myVec_57 : _GEN_1570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1572 = 6'h3a == _myNewVec_41_T_3[5:0] ? myVec_58 : _GEN_1571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1573 = 6'h3b == _myNewVec_41_T_3[5:0] ? myVec_59 : _GEN_1572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1574 = 6'h3c == _myNewVec_41_T_3[5:0] ? myVec_60 : _GEN_1573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1575 = 6'h3d == _myNewVec_41_T_3[5:0] ? myVec_61 : _GEN_1574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1576 = 6'h3e == _myNewVec_41_T_3[5:0] ? myVec_62 : _GEN_1575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_41 = 6'h3f == _myNewVec_41_T_3[5:0] ? myVec_63 : _GEN_1576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_40_T_3 = _myNewVec_63_T_1 + 16'h17; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1579 = 6'h1 == _myNewVec_40_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1580 = 6'h2 == _myNewVec_40_T_3[5:0] ? myVec_2 : _GEN_1579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1581 = 6'h3 == _myNewVec_40_T_3[5:0] ? myVec_3 : _GEN_1580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1582 = 6'h4 == _myNewVec_40_T_3[5:0] ? myVec_4 : _GEN_1581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1583 = 6'h5 == _myNewVec_40_T_3[5:0] ? myVec_5 : _GEN_1582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1584 = 6'h6 == _myNewVec_40_T_3[5:0] ? myVec_6 : _GEN_1583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1585 = 6'h7 == _myNewVec_40_T_3[5:0] ? myVec_7 : _GEN_1584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1586 = 6'h8 == _myNewVec_40_T_3[5:0] ? myVec_8 : _GEN_1585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1587 = 6'h9 == _myNewVec_40_T_3[5:0] ? myVec_9 : _GEN_1586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1588 = 6'ha == _myNewVec_40_T_3[5:0] ? myVec_10 : _GEN_1587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1589 = 6'hb == _myNewVec_40_T_3[5:0] ? myVec_11 : _GEN_1588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1590 = 6'hc == _myNewVec_40_T_3[5:0] ? myVec_12 : _GEN_1589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1591 = 6'hd == _myNewVec_40_T_3[5:0] ? myVec_13 : _GEN_1590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1592 = 6'he == _myNewVec_40_T_3[5:0] ? myVec_14 : _GEN_1591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1593 = 6'hf == _myNewVec_40_T_3[5:0] ? myVec_15 : _GEN_1592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1594 = 6'h10 == _myNewVec_40_T_3[5:0] ? myVec_16 : _GEN_1593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1595 = 6'h11 == _myNewVec_40_T_3[5:0] ? myVec_17 : _GEN_1594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1596 = 6'h12 == _myNewVec_40_T_3[5:0] ? myVec_18 : _GEN_1595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1597 = 6'h13 == _myNewVec_40_T_3[5:0] ? myVec_19 : _GEN_1596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1598 = 6'h14 == _myNewVec_40_T_3[5:0] ? myVec_20 : _GEN_1597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1599 = 6'h15 == _myNewVec_40_T_3[5:0] ? myVec_21 : _GEN_1598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1600 = 6'h16 == _myNewVec_40_T_3[5:0] ? myVec_22 : _GEN_1599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1601 = 6'h17 == _myNewVec_40_T_3[5:0] ? myVec_23 : _GEN_1600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1602 = 6'h18 == _myNewVec_40_T_3[5:0] ? myVec_24 : _GEN_1601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1603 = 6'h19 == _myNewVec_40_T_3[5:0] ? myVec_25 : _GEN_1602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1604 = 6'h1a == _myNewVec_40_T_3[5:0] ? myVec_26 : _GEN_1603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1605 = 6'h1b == _myNewVec_40_T_3[5:0] ? myVec_27 : _GEN_1604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1606 = 6'h1c == _myNewVec_40_T_3[5:0] ? myVec_28 : _GEN_1605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1607 = 6'h1d == _myNewVec_40_T_3[5:0] ? myVec_29 : _GEN_1606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1608 = 6'h1e == _myNewVec_40_T_3[5:0] ? myVec_30 : _GEN_1607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1609 = 6'h1f == _myNewVec_40_T_3[5:0] ? myVec_31 : _GEN_1608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1610 = 6'h20 == _myNewVec_40_T_3[5:0] ? myVec_32 : _GEN_1609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1611 = 6'h21 == _myNewVec_40_T_3[5:0] ? myVec_33 : _GEN_1610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1612 = 6'h22 == _myNewVec_40_T_3[5:0] ? myVec_34 : _GEN_1611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1613 = 6'h23 == _myNewVec_40_T_3[5:0] ? myVec_35 : _GEN_1612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1614 = 6'h24 == _myNewVec_40_T_3[5:0] ? myVec_36 : _GEN_1613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1615 = 6'h25 == _myNewVec_40_T_3[5:0] ? myVec_37 : _GEN_1614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1616 = 6'h26 == _myNewVec_40_T_3[5:0] ? myVec_38 : _GEN_1615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1617 = 6'h27 == _myNewVec_40_T_3[5:0] ? myVec_39 : _GEN_1616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1618 = 6'h28 == _myNewVec_40_T_3[5:0] ? myVec_40 : _GEN_1617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1619 = 6'h29 == _myNewVec_40_T_3[5:0] ? myVec_41 : _GEN_1618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1620 = 6'h2a == _myNewVec_40_T_3[5:0] ? myVec_42 : _GEN_1619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1621 = 6'h2b == _myNewVec_40_T_3[5:0] ? myVec_43 : _GEN_1620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1622 = 6'h2c == _myNewVec_40_T_3[5:0] ? myVec_44 : _GEN_1621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1623 = 6'h2d == _myNewVec_40_T_3[5:0] ? myVec_45 : _GEN_1622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1624 = 6'h2e == _myNewVec_40_T_3[5:0] ? myVec_46 : _GEN_1623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1625 = 6'h2f == _myNewVec_40_T_3[5:0] ? myVec_47 : _GEN_1624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1626 = 6'h30 == _myNewVec_40_T_3[5:0] ? myVec_48 : _GEN_1625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1627 = 6'h31 == _myNewVec_40_T_3[5:0] ? myVec_49 : _GEN_1626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1628 = 6'h32 == _myNewVec_40_T_3[5:0] ? myVec_50 : _GEN_1627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1629 = 6'h33 == _myNewVec_40_T_3[5:0] ? myVec_51 : _GEN_1628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1630 = 6'h34 == _myNewVec_40_T_3[5:0] ? myVec_52 : _GEN_1629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1631 = 6'h35 == _myNewVec_40_T_3[5:0] ? myVec_53 : _GEN_1630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1632 = 6'h36 == _myNewVec_40_T_3[5:0] ? myVec_54 : _GEN_1631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1633 = 6'h37 == _myNewVec_40_T_3[5:0] ? myVec_55 : _GEN_1632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1634 = 6'h38 == _myNewVec_40_T_3[5:0] ? myVec_56 : _GEN_1633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1635 = 6'h39 == _myNewVec_40_T_3[5:0] ? myVec_57 : _GEN_1634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1636 = 6'h3a == _myNewVec_40_T_3[5:0] ? myVec_58 : _GEN_1635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1637 = 6'h3b == _myNewVec_40_T_3[5:0] ? myVec_59 : _GEN_1636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1638 = 6'h3c == _myNewVec_40_T_3[5:0] ? myVec_60 : _GEN_1637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1639 = 6'h3d == _myNewVec_40_T_3[5:0] ? myVec_61 : _GEN_1638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1640 = 6'h3e == _myNewVec_40_T_3[5:0] ? myVec_62 : _GEN_1639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_40 = 6'h3f == _myNewVec_40_T_3[5:0] ? myVec_63 : _GEN_1640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_39_T_3 = _myNewVec_63_T_1 + 16'h18; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1643 = 6'h1 == _myNewVec_39_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1644 = 6'h2 == _myNewVec_39_T_3[5:0] ? myVec_2 : _GEN_1643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1645 = 6'h3 == _myNewVec_39_T_3[5:0] ? myVec_3 : _GEN_1644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1646 = 6'h4 == _myNewVec_39_T_3[5:0] ? myVec_4 : _GEN_1645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1647 = 6'h5 == _myNewVec_39_T_3[5:0] ? myVec_5 : _GEN_1646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1648 = 6'h6 == _myNewVec_39_T_3[5:0] ? myVec_6 : _GEN_1647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1649 = 6'h7 == _myNewVec_39_T_3[5:0] ? myVec_7 : _GEN_1648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1650 = 6'h8 == _myNewVec_39_T_3[5:0] ? myVec_8 : _GEN_1649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1651 = 6'h9 == _myNewVec_39_T_3[5:0] ? myVec_9 : _GEN_1650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1652 = 6'ha == _myNewVec_39_T_3[5:0] ? myVec_10 : _GEN_1651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1653 = 6'hb == _myNewVec_39_T_3[5:0] ? myVec_11 : _GEN_1652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1654 = 6'hc == _myNewVec_39_T_3[5:0] ? myVec_12 : _GEN_1653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1655 = 6'hd == _myNewVec_39_T_3[5:0] ? myVec_13 : _GEN_1654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1656 = 6'he == _myNewVec_39_T_3[5:0] ? myVec_14 : _GEN_1655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1657 = 6'hf == _myNewVec_39_T_3[5:0] ? myVec_15 : _GEN_1656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1658 = 6'h10 == _myNewVec_39_T_3[5:0] ? myVec_16 : _GEN_1657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1659 = 6'h11 == _myNewVec_39_T_3[5:0] ? myVec_17 : _GEN_1658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1660 = 6'h12 == _myNewVec_39_T_3[5:0] ? myVec_18 : _GEN_1659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1661 = 6'h13 == _myNewVec_39_T_3[5:0] ? myVec_19 : _GEN_1660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1662 = 6'h14 == _myNewVec_39_T_3[5:0] ? myVec_20 : _GEN_1661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1663 = 6'h15 == _myNewVec_39_T_3[5:0] ? myVec_21 : _GEN_1662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1664 = 6'h16 == _myNewVec_39_T_3[5:0] ? myVec_22 : _GEN_1663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1665 = 6'h17 == _myNewVec_39_T_3[5:0] ? myVec_23 : _GEN_1664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1666 = 6'h18 == _myNewVec_39_T_3[5:0] ? myVec_24 : _GEN_1665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1667 = 6'h19 == _myNewVec_39_T_3[5:0] ? myVec_25 : _GEN_1666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1668 = 6'h1a == _myNewVec_39_T_3[5:0] ? myVec_26 : _GEN_1667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1669 = 6'h1b == _myNewVec_39_T_3[5:0] ? myVec_27 : _GEN_1668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1670 = 6'h1c == _myNewVec_39_T_3[5:0] ? myVec_28 : _GEN_1669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1671 = 6'h1d == _myNewVec_39_T_3[5:0] ? myVec_29 : _GEN_1670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1672 = 6'h1e == _myNewVec_39_T_3[5:0] ? myVec_30 : _GEN_1671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1673 = 6'h1f == _myNewVec_39_T_3[5:0] ? myVec_31 : _GEN_1672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1674 = 6'h20 == _myNewVec_39_T_3[5:0] ? myVec_32 : _GEN_1673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1675 = 6'h21 == _myNewVec_39_T_3[5:0] ? myVec_33 : _GEN_1674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1676 = 6'h22 == _myNewVec_39_T_3[5:0] ? myVec_34 : _GEN_1675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1677 = 6'h23 == _myNewVec_39_T_3[5:0] ? myVec_35 : _GEN_1676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1678 = 6'h24 == _myNewVec_39_T_3[5:0] ? myVec_36 : _GEN_1677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1679 = 6'h25 == _myNewVec_39_T_3[5:0] ? myVec_37 : _GEN_1678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1680 = 6'h26 == _myNewVec_39_T_3[5:0] ? myVec_38 : _GEN_1679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1681 = 6'h27 == _myNewVec_39_T_3[5:0] ? myVec_39 : _GEN_1680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1682 = 6'h28 == _myNewVec_39_T_3[5:0] ? myVec_40 : _GEN_1681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1683 = 6'h29 == _myNewVec_39_T_3[5:0] ? myVec_41 : _GEN_1682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1684 = 6'h2a == _myNewVec_39_T_3[5:0] ? myVec_42 : _GEN_1683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1685 = 6'h2b == _myNewVec_39_T_3[5:0] ? myVec_43 : _GEN_1684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1686 = 6'h2c == _myNewVec_39_T_3[5:0] ? myVec_44 : _GEN_1685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1687 = 6'h2d == _myNewVec_39_T_3[5:0] ? myVec_45 : _GEN_1686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1688 = 6'h2e == _myNewVec_39_T_3[5:0] ? myVec_46 : _GEN_1687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1689 = 6'h2f == _myNewVec_39_T_3[5:0] ? myVec_47 : _GEN_1688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1690 = 6'h30 == _myNewVec_39_T_3[5:0] ? myVec_48 : _GEN_1689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1691 = 6'h31 == _myNewVec_39_T_3[5:0] ? myVec_49 : _GEN_1690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1692 = 6'h32 == _myNewVec_39_T_3[5:0] ? myVec_50 : _GEN_1691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1693 = 6'h33 == _myNewVec_39_T_3[5:0] ? myVec_51 : _GEN_1692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1694 = 6'h34 == _myNewVec_39_T_3[5:0] ? myVec_52 : _GEN_1693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1695 = 6'h35 == _myNewVec_39_T_3[5:0] ? myVec_53 : _GEN_1694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1696 = 6'h36 == _myNewVec_39_T_3[5:0] ? myVec_54 : _GEN_1695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1697 = 6'h37 == _myNewVec_39_T_3[5:0] ? myVec_55 : _GEN_1696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1698 = 6'h38 == _myNewVec_39_T_3[5:0] ? myVec_56 : _GEN_1697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1699 = 6'h39 == _myNewVec_39_T_3[5:0] ? myVec_57 : _GEN_1698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1700 = 6'h3a == _myNewVec_39_T_3[5:0] ? myVec_58 : _GEN_1699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1701 = 6'h3b == _myNewVec_39_T_3[5:0] ? myVec_59 : _GEN_1700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1702 = 6'h3c == _myNewVec_39_T_3[5:0] ? myVec_60 : _GEN_1701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1703 = 6'h3d == _myNewVec_39_T_3[5:0] ? myVec_61 : _GEN_1702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1704 = 6'h3e == _myNewVec_39_T_3[5:0] ? myVec_62 : _GEN_1703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_39 = 6'h3f == _myNewVec_39_T_3[5:0] ? myVec_63 : _GEN_1704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_38_T_3 = _myNewVec_63_T_1 + 16'h19; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1707 = 6'h1 == _myNewVec_38_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1708 = 6'h2 == _myNewVec_38_T_3[5:0] ? myVec_2 : _GEN_1707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1709 = 6'h3 == _myNewVec_38_T_3[5:0] ? myVec_3 : _GEN_1708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1710 = 6'h4 == _myNewVec_38_T_3[5:0] ? myVec_4 : _GEN_1709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1711 = 6'h5 == _myNewVec_38_T_3[5:0] ? myVec_5 : _GEN_1710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1712 = 6'h6 == _myNewVec_38_T_3[5:0] ? myVec_6 : _GEN_1711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1713 = 6'h7 == _myNewVec_38_T_3[5:0] ? myVec_7 : _GEN_1712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1714 = 6'h8 == _myNewVec_38_T_3[5:0] ? myVec_8 : _GEN_1713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1715 = 6'h9 == _myNewVec_38_T_3[5:0] ? myVec_9 : _GEN_1714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1716 = 6'ha == _myNewVec_38_T_3[5:0] ? myVec_10 : _GEN_1715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1717 = 6'hb == _myNewVec_38_T_3[5:0] ? myVec_11 : _GEN_1716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1718 = 6'hc == _myNewVec_38_T_3[5:0] ? myVec_12 : _GEN_1717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1719 = 6'hd == _myNewVec_38_T_3[5:0] ? myVec_13 : _GEN_1718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1720 = 6'he == _myNewVec_38_T_3[5:0] ? myVec_14 : _GEN_1719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1721 = 6'hf == _myNewVec_38_T_3[5:0] ? myVec_15 : _GEN_1720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1722 = 6'h10 == _myNewVec_38_T_3[5:0] ? myVec_16 : _GEN_1721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1723 = 6'h11 == _myNewVec_38_T_3[5:0] ? myVec_17 : _GEN_1722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1724 = 6'h12 == _myNewVec_38_T_3[5:0] ? myVec_18 : _GEN_1723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1725 = 6'h13 == _myNewVec_38_T_3[5:0] ? myVec_19 : _GEN_1724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1726 = 6'h14 == _myNewVec_38_T_3[5:0] ? myVec_20 : _GEN_1725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1727 = 6'h15 == _myNewVec_38_T_3[5:0] ? myVec_21 : _GEN_1726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1728 = 6'h16 == _myNewVec_38_T_3[5:0] ? myVec_22 : _GEN_1727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1729 = 6'h17 == _myNewVec_38_T_3[5:0] ? myVec_23 : _GEN_1728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1730 = 6'h18 == _myNewVec_38_T_3[5:0] ? myVec_24 : _GEN_1729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1731 = 6'h19 == _myNewVec_38_T_3[5:0] ? myVec_25 : _GEN_1730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1732 = 6'h1a == _myNewVec_38_T_3[5:0] ? myVec_26 : _GEN_1731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1733 = 6'h1b == _myNewVec_38_T_3[5:0] ? myVec_27 : _GEN_1732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1734 = 6'h1c == _myNewVec_38_T_3[5:0] ? myVec_28 : _GEN_1733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1735 = 6'h1d == _myNewVec_38_T_3[5:0] ? myVec_29 : _GEN_1734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1736 = 6'h1e == _myNewVec_38_T_3[5:0] ? myVec_30 : _GEN_1735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1737 = 6'h1f == _myNewVec_38_T_3[5:0] ? myVec_31 : _GEN_1736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1738 = 6'h20 == _myNewVec_38_T_3[5:0] ? myVec_32 : _GEN_1737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1739 = 6'h21 == _myNewVec_38_T_3[5:0] ? myVec_33 : _GEN_1738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1740 = 6'h22 == _myNewVec_38_T_3[5:0] ? myVec_34 : _GEN_1739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1741 = 6'h23 == _myNewVec_38_T_3[5:0] ? myVec_35 : _GEN_1740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1742 = 6'h24 == _myNewVec_38_T_3[5:0] ? myVec_36 : _GEN_1741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1743 = 6'h25 == _myNewVec_38_T_3[5:0] ? myVec_37 : _GEN_1742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1744 = 6'h26 == _myNewVec_38_T_3[5:0] ? myVec_38 : _GEN_1743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1745 = 6'h27 == _myNewVec_38_T_3[5:0] ? myVec_39 : _GEN_1744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1746 = 6'h28 == _myNewVec_38_T_3[5:0] ? myVec_40 : _GEN_1745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1747 = 6'h29 == _myNewVec_38_T_3[5:0] ? myVec_41 : _GEN_1746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1748 = 6'h2a == _myNewVec_38_T_3[5:0] ? myVec_42 : _GEN_1747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1749 = 6'h2b == _myNewVec_38_T_3[5:0] ? myVec_43 : _GEN_1748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1750 = 6'h2c == _myNewVec_38_T_3[5:0] ? myVec_44 : _GEN_1749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1751 = 6'h2d == _myNewVec_38_T_3[5:0] ? myVec_45 : _GEN_1750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1752 = 6'h2e == _myNewVec_38_T_3[5:0] ? myVec_46 : _GEN_1751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1753 = 6'h2f == _myNewVec_38_T_3[5:0] ? myVec_47 : _GEN_1752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1754 = 6'h30 == _myNewVec_38_T_3[5:0] ? myVec_48 : _GEN_1753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1755 = 6'h31 == _myNewVec_38_T_3[5:0] ? myVec_49 : _GEN_1754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1756 = 6'h32 == _myNewVec_38_T_3[5:0] ? myVec_50 : _GEN_1755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1757 = 6'h33 == _myNewVec_38_T_3[5:0] ? myVec_51 : _GEN_1756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1758 = 6'h34 == _myNewVec_38_T_3[5:0] ? myVec_52 : _GEN_1757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1759 = 6'h35 == _myNewVec_38_T_3[5:0] ? myVec_53 : _GEN_1758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1760 = 6'h36 == _myNewVec_38_T_3[5:0] ? myVec_54 : _GEN_1759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1761 = 6'h37 == _myNewVec_38_T_3[5:0] ? myVec_55 : _GEN_1760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1762 = 6'h38 == _myNewVec_38_T_3[5:0] ? myVec_56 : _GEN_1761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1763 = 6'h39 == _myNewVec_38_T_3[5:0] ? myVec_57 : _GEN_1762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1764 = 6'h3a == _myNewVec_38_T_3[5:0] ? myVec_58 : _GEN_1763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1765 = 6'h3b == _myNewVec_38_T_3[5:0] ? myVec_59 : _GEN_1764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1766 = 6'h3c == _myNewVec_38_T_3[5:0] ? myVec_60 : _GEN_1765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1767 = 6'h3d == _myNewVec_38_T_3[5:0] ? myVec_61 : _GEN_1766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1768 = 6'h3e == _myNewVec_38_T_3[5:0] ? myVec_62 : _GEN_1767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_38 = 6'h3f == _myNewVec_38_T_3[5:0] ? myVec_63 : _GEN_1768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_37_T_3 = _myNewVec_63_T_1 + 16'h1a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1771 = 6'h1 == _myNewVec_37_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1772 = 6'h2 == _myNewVec_37_T_3[5:0] ? myVec_2 : _GEN_1771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1773 = 6'h3 == _myNewVec_37_T_3[5:0] ? myVec_3 : _GEN_1772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1774 = 6'h4 == _myNewVec_37_T_3[5:0] ? myVec_4 : _GEN_1773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1775 = 6'h5 == _myNewVec_37_T_3[5:0] ? myVec_5 : _GEN_1774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1776 = 6'h6 == _myNewVec_37_T_3[5:0] ? myVec_6 : _GEN_1775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1777 = 6'h7 == _myNewVec_37_T_3[5:0] ? myVec_7 : _GEN_1776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1778 = 6'h8 == _myNewVec_37_T_3[5:0] ? myVec_8 : _GEN_1777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1779 = 6'h9 == _myNewVec_37_T_3[5:0] ? myVec_9 : _GEN_1778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1780 = 6'ha == _myNewVec_37_T_3[5:0] ? myVec_10 : _GEN_1779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1781 = 6'hb == _myNewVec_37_T_3[5:0] ? myVec_11 : _GEN_1780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1782 = 6'hc == _myNewVec_37_T_3[5:0] ? myVec_12 : _GEN_1781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1783 = 6'hd == _myNewVec_37_T_3[5:0] ? myVec_13 : _GEN_1782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1784 = 6'he == _myNewVec_37_T_3[5:0] ? myVec_14 : _GEN_1783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1785 = 6'hf == _myNewVec_37_T_3[5:0] ? myVec_15 : _GEN_1784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1786 = 6'h10 == _myNewVec_37_T_3[5:0] ? myVec_16 : _GEN_1785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1787 = 6'h11 == _myNewVec_37_T_3[5:0] ? myVec_17 : _GEN_1786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1788 = 6'h12 == _myNewVec_37_T_3[5:0] ? myVec_18 : _GEN_1787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1789 = 6'h13 == _myNewVec_37_T_3[5:0] ? myVec_19 : _GEN_1788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1790 = 6'h14 == _myNewVec_37_T_3[5:0] ? myVec_20 : _GEN_1789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1791 = 6'h15 == _myNewVec_37_T_3[5:0] ? myVec_21 : _GEN_1790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1792 = 6'h16 == _myNewVec_37_T_3[5:0] ? myVec_22 : _GEN_1791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1793 = 6'h17 == _myNewVec_37_T_3[5:0] ? myVec_23 : _GEN_1792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1794 = 6'h18 == _myNewVec_37_T_3[5:0] ? myVec_24 : _GEN_1793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1795 = 6'h19 == _myNewVec_37_T_3[5:0] ? myVec_25 : _GEN_1794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1796 = 6'h1a == _myNewVec_37_T_3[5:0] ? myVec_26 : _GEN_1795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1797 = 6'h1b == _myNewVec_37_T_3[5:0] ? myVec_27 : _GEN_1796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1798 = 6'h1c == _myNewVec_37_T_3[5:0] ? myVec_28 : _GEN_1797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1799 = 6'h1d == _myNewVec_37_T_3[5:0] ? myVec_29 : _GEN_1798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1800 = 6'h1e == _myNewVec_37_T_3[5:0] ? myVec_30 : _GEN_1799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1801 = 6'h1f == _myNewVec_37_T_3[5:0] ? myVec_31 : _GEN_1800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1802 = 6'h20 == _myNewVec_37_T_3[5:0] ? myVec_32 : _GEN_1801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1803 = 6'h21 == _myNewVec_37_T_3[5:0] ? myVec_33 : _GEN_1802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1804 = 6'h22 == _myNewVec_37_T_3[5:0] ? myVec_34 : _GEN_1803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1805 = 6'h23 == _myNewVec_37_T_3[5:0] ? myVec_35 : _GEN_1804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1806 = 6'h24 == _myNewVec_37_T_3[5:0] ? myVec_36 : _GEN_1805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1807 = 6'h25 == _myNewVec_37_T_3[5:0] ? myVec_37 : _GEN_1806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1808 = 6'h26 == _myNewVec_37_T_3[5:0] ? myVec_38 : _GEN_1807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1809 = 6'h27 == _myNewVec_37_T_3[5:0] ? myVec_39 : _GEN_1808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1810 = 6'h28 == _myNewVec_37_T_3[5:0] ? myVec_40 : _GEN_1809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1811 = 6'h29 == _myNewVec_37_T_3[5:0] ? myVec_41 : _GEN_1810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1812 = 6'h2a == _myNewVec_37_T_3[5:0] ? myVec_42 : _GEN_1811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1813 = 6'h2b == _myNewVec_37_T_3[5:0] ? myVec_43 : _GEN_1812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1814 = 6'h2c == _myNewVec_37_T_3[5:0] ? myVec_44 : _GEN_1813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1815 = 6'h2d == _myNewVec_37_T_3[5:0] ? myVec_45 : _GEN_1814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1816 = 6'h2e == _myNewVec_37_T_3[5:0] ? myVec_46 : _GEN_1815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1817 = 6'h2f == _myNewVec_37_T_3[5:0] ? myVec_47 : _GEN_1816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1818 = 6'h30 == _myNewVec_37_T_3[5:0] ? myVec_48 : _GEN_1817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1819 = 6'h31 == _myNewVec_37_T_3[5:0] ? myVec_49 : _GEN_1818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1820 = 6'h32 == _myNewVec_37_T_3[5:0] ? myVec_50 : _GEN_1819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1821 = 6'h33 == _myNewVec_37_T_3[5:0] ? myVec_51 : _GEN_1820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1822 = 6'h34 == _myNewVec_37_T_3[5:0] ? myVec_52 : _GEN_1821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1823 = 6'h35 == _myNewVec_37_T_3[5:0] ? myVec_53 : _GEN_1822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1824 = 6'h36 == _myNewVec_37_T_3[5:0] ? myVec_54 : _GEN_1823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1825 = 6'h37 == _myNewVec_37_T_3[5:0] ? myVec_55 : _GEN_1824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1826 = 6'h38 == _myNewVec_37_T_3[5:0] ? myVec_56 : _GEN_1825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1827 = 6'h39 == _myNewVec_37_T_3[5:0] ? myVec_57 : _GEN_1826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1828 = 6'h3a == _myNewVec_37_T_3[5:0] ? myVec_58 : _GEN_1827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1829 = 6'h3b == _myNewVec_37_T_3[5:0] ? myVec_59 : _GEN_1828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1830 = 6'h3c == _myNewVec_37_T_3[5:0] ? myVec_60 : _GEN_1829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1831 = 6'h3d == _myNewVec_37_T_3[5:0] ? myVec_61 : _GEN_1830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1832 = 6'h3e == _myNewVec_37_T_3[5:0] ? myVec_62 : _GEN_1831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_37 = 6'h3f == _myNewVec_37_T_3[5:0] ? myVec_63 : _GEN_1832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_36_T_3 = _myNewVec_63_T_1 + 16'h1b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1835 = 6'h1 == _myNewVec_36_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1836 = 6'h2 == _myNewVec_36_T_3[5:0] ? myVec_2 : _GEN_1835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1837 = 6'h3 == _myNewVec_36_T_3[5:0] ? myVec_3 : _GEN_1836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1838 = 6'h4 == _myNewVec_36_T_3[5:0] ? myVec_4 : _GEN_1837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1839 = 6'h5 == _myNewVec_36_T_3[5:0] ? myVec_5 : _GEN_1838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1840 = 6'h6 == _myNewVec_36_T_3[5:0] ? myVec_6 : _GEN_1839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1841 = 6'h7 == _myNewVec_36_T_3[5:0] ? myVec_7 : _GEN_1840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1842 = 6'h8 == _myNewVec_36_T_3[5:0] ? myVec_8 : _GEN_1841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1843 = 6'h9 == _myNewVec_36_T_3[5:0] ? myVec_9 : _GEN_1842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1844 = 6'ha == _myNewVec_36_T_3[5:0] ? myVec_10 : _GEN_1843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1845 = 6'hb == _myNewVec_36_T_3[5:0] ? myVec_11 : _GEN_1844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1846 = 6'hc == _myNewVec_36_T_3[5:0] ? myVec_12 : _GEN_1845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1847 = 6'hd == _myNewVec_36_T_3[5:0] ? myVec_13 : _GEN_1846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1848 = 6'he == _myNewVec_36_T_3[5:0] ? myVec_14 : _GEN_1847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1849 = 6'hf == _myNewVec_36_T_3[5:0] ? myVec_15 : _GEN_1848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1850 = 6'h10 == _myNewVec_36_T_3[5:0] ? myVec_16 : _GEN_1849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1851 = 6'h11 == _myNewVec_36_T_3[5:0] ? myVec_17 : _GEN_1850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1852 = 6'h12 == _myNewVec_36_T_3[5:0] ? myVec_18 : _GEN_1851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1853 = 6'h13 == _myNewVec_36_T_3[5:0] ? myVec_19 : _GEN_1852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1854 = 6'h14 == _myNewVec_36_T_3[5:0] ? myVec_20 : _GEN_1853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1855 = 6'h15 == _myNewVec_36_T_3[5:0] ? myVec_21 : _GEN_1854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1856 = 6'h16 == _myNewVec_36_T_3[5:0] ? myVec_22 : _GEN_1855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1857 = 6'h17 == _myNewVec_36_T_3[5:0] ? myVec_23 : _GEN_1856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1858 = 6'h18 == _myNewVec_36_T_3[5:0] ? myVec_24 : _GEN_1857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1859 = 6'h19 == _myNewVec_36_T_3[5:0] ? myVec_25 : _GEN_1858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1860 = 6'h1a == _myNewVec_36_T_3[5:0] ? myVec_26 : _GEN_1859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1861 = 6'h1b == _myNewVec_36_T_3[5:0] ? myVec_27 : _GEN_1860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1862 = 6'h1c == _myNewVec_36_T_3[5:0] ? myVec_28 : _GEN_1861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1863 = 6'h1d == _myNewVec_36_T_3[5:0] ? myVec_29 : _GEN_1862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1864 = 6'h1e == _myNewVec_36_T_3[5:0] ? myVec_30 : _GEN_1863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1865 = 6'h1f == _myNewVec_36_T_3[5:0] ? myVec_31 : _GEN_1864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1866 = 6'h20 == _myNewVec_36_T_3[5:0] ? myVec_32 : _GEN_1865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1867 = 6'h21 == _myNewVec_36_T_3[5:0] ? myVec_33 : _GEN_1866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1868 = 6'h22 == _myNewVec_36_T_3[5:0] ? myVec_34 : _GEN_1867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1869 = 6'h23 == _myNewVec_36_T_3[5:0] ? myVec_35 : _GEN_1868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1870 = 6'h24 == _myNewVec_36_T_3[5:0] ? myVec_36 : _GEN_1869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1871 = 6'h25 == _myNewVec_36_T_3[5:0] ? myVec_37 : _GEN_1870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1872 = 6'h26 == _myNewVec_36_T_3[5:0] ? myVec_38 : _GEN_1871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1873 = 6'h27 == _myNewVec_36_T_3[5:0] ? myVec_39 : _GEN_1872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1874 = 6'h28 == _myNewVec_36_T_3[5:0] ? myVec_40 : _GEN_1873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1875 = 6'h29 == _myNewVec_36_T_3[5:0] ? myVec_41 : _GEN_1874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1876 = 6'h2a == _myNewVec_36_T_3[5:0] ? myVec_42 : _GEN_1875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1877 = 6'h2b == _myNewVec_36_T_3[5:0] ? myVec_43 : _GEN_1876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1878 = 6'h2c == _myNewVec_36_T_3[5:0] ? myVec_44 : _GEN_1877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1879 = 6'h2d == _myNewVec_36_T_3[5:0] ? myVec_45 : _GEN_1878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1880 = 6'h2e == _myNewVec_36_T_3[5:0] ? myVec_46 : _GEN_1879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1881 = 6'h2f == _myNewVec_36_T_3[5:0] ? myVec_47 : _GEN_1880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1882 = 6'h30 == _myNewVec_36_T_3[5:0] ? myVec_48 : _GEN_1881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1883 = 6'h31 == _myNewVec_36_T_3[5:0] ? myVec_49 : _GEN_1882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1884 = 6'h32 == _myNewVec_36_T_3[5:0] ? myVec_50 : _GEN_1883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1885 = 6'h33 == _myNewVec_36_T_3[5:0] ? myVec_51 : _GEN_1884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1886 = 6'h34 == _myNewVec_36_T_3[5:0] ? myVec_52 : _GEN_1885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1887 = 6'h35 == _myNewVec_36_T_3[5:0] ? myVec_53 : _GEN_1886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1888 = 6'h36 == _myNewVec_36_T_3[5:0] ? myVec_54 : _GEN_1887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1889 = 6'h37 == _myNewVec_36_T_3[5:0] ? myVec_55 : _GEN_1888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1890 = 6'h38 == _myNewVec_36_T_3[5:0] ? myVec_56 : _GEN_1889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1891 = 6'h39 == _myNewVec_36_T_3[5:0] ? myVec_57 : _GEN_1890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1892 = 6'h3a == _myNewVec_36_T_3[5:0] ? myVec_58 : _GEN_1891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1893 = 6'h3b == _myNewVec_36_T_3[5:0] ? myVec_59 : _GEN_1892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1894 = 6'h3c == _myNewVec_36_T_3[5:0] ? myVec_60 : _GEN_1893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1895 = 6'h3d == _myNewVec_36_T_3[5:0] ? myVec_61 : _GEN_1894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1896 = 6'h3e == _myNewVec_36_T_3[5:0] ? myVec_62 : _GEN_1895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_36 = 6'h3f == _myNewVec_36_T_3[5:0] ? myVec_63 : _GEN_1896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_35_T_3 = _myNewVec_63_T_1 + 16'h1c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1899 = 6'h1 == _myNewVec_35_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1900 = 6'h2 == _myNewVec_35_T_3[5:0] ? myVec_2 : _GEN_1899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1901 = 6'h3 == _myNewVec_35_T_3[5:0] ? myVec_3 : _GEN_1900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1902 = 6'h4 == _myNewVec_35_T_3[5:0] ? myVec_4 : _GEN_1901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1903 = 6'h5 == _myNewVec_35_T_3[5:0] ? myVec_5 : _GEN_1902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1904 = 6'h6 == _myNewVec_35_T_3[5:0] ? myVec_6 : _GEN_1903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1905 = 6'h7 == _myNewVec_35_T_3[5:0] ? myVec_7 : _GEN_1904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1906 = 6'h8 == _myNewVec_35_T_3[5:0] ? myVec_8 : _GEN_1905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1907 = 6'h9 == _myNewVec_35_T_3[5:0] ? myVec_9 : _GEN_1906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1908 = 6'ha == _myNewVec_35_T_3[5:0] ? myVec_10 : _GEN_1907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1909 = 6'hb == _myNewVec_35_T_3[5:0] ? myVec_11 : _GEN_1908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1910 = 6'hc == _myNewVec_35_T_3[5:0] ? myVec_12 : _GEN_1909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1911 = 6'hd == _myNewVec_35_T_3[5:0] ? myVec_13 : _GEN_1910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1912 = 6'he == _myNewVec_35_T_3[5:0] ? myVec_14 : _GEN_1911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1913 = 6'hf == _myNewVec_35_T_3[5:0] ? myVec_15 : _GEN_1912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1914 = 6'h10 == _myNewVec_35_T_3[5:0] ? myVec_16 : _GEN_1913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1915 = 6'h11 == _myNewVec_35_T_3[5:0] ? myVec_17 : _GEN_1914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1916 = 6'h12 == _myNewVec_35_T_3[5:0] ? myVec_18 : _GEN_1915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1917 = 6'h13 == _myNewVec_35_T_3[5:0] ? myVec_19 : _GEN_1916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1918 = 6'h14 == _myNewVec_35_T_3[5:0] ? myVec_20 : _GEN_1917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1919 = 6'h15 == _myNewVec_35_T_3[5:0] ? myVec_21 : _GEN_1918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1920 = 6'h16 == _myNewVec_35_T_3[5:0] ? myVec_22 : _GEN_1919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1921 = 6'h17 == _myNewVec_35_T_3[5:0] ? myVec_23 : _GEN_1920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1922 = 6'h18 == _myNewVec_35_T_3[5:0] ? myVec_24 : _GEN_1921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1923 = 6'h19 == _myNewVec_35_T_3[5:0] ? myVec_25 : _GEN_1922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1924 = 6'h1a == _myNewVec_35_T_3[5:0] ? myVec_26 : _GEN_1923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1925 = 6'h1b == _myNewVec_35_T_3[5:0] ? myVec_27 : _GEN_1924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1926 = 6'h1c == _myNewVec_35_T_3[5:0] ? myVec_28 : _GEN_1925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1927 = 6'h1d == _myNewVec_35_T_3[5:0] ? myVec_29 : _GEN_1926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1928 = 6'h1e == _myNewVec_35_T_3[5:0] ? myVec_30 : _GEN_1927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1929 = 6'h1f == _myNewVec_35_T_3[5:0] ? myVec_31 : _GEN_1928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1930 = 6'h20 == _myNewVec_35_T_3[5:0] ? myVec_32 : _GEN_1929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1931 = 6'h21 == _myNewVec_35_T_3[5:0] ? myVec_33 : _GEN_1930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1932 = 6'h22 == _myNewVec_35_T_3[5:0] ? myVec_34 : _GEN_1931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1933 = 6'h23 == _myNewVec_35_T_3[5:0] ? myVec_35 : _GEN_1932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1934 = 6'h24 == _myNewVec_35_T_3[5:0] ? myVec_36 : _GEN_1933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1935 = 6'h25 == _myNewVec_35_T_3[5:0] ? myVec_37 : _GEN_1934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1936 = 6'h26 == _myNewVec_35_T_3[5:0] ? myVec_38 : _GEN_1935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1937 = 6'h27 == _myNewVec_35_T_3[5:0] ? myVec_39 : _GEN_1936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1938 = 6'h28 == _myNewVec_35_T_3[5:0] ? myVec_40 : _GEN_1937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1939 = 6'h29 == _myNewVec_35_T_3[5:0] ? myVec_41 : _GEN_1938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1940 = 6'h2a == _myNewVec_35_T_3[5:0] ? myVec_42 : _GEN_1939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1941 = 6'h2b == _myNewVec_35_T_3[5:0] ? myVec_43 : _GEN_1940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1942 = 6'h2c == _myNewVec_35_T_3[5:0] ? myVec_44 : _GEN_1941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1943 = 6'h2d == _myNewVec_35_T_3[5:0] ? myVec_45 : _GEN_1942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1944 = 6'h2e == _myNewVec_35_T_3[5:0] ? myVec_46 : _GEN_1943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1945 = 6'h2f == _myNewVec_35_T_3[5:0] ? myVec_47 : _GEN_1944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1946 = 6'h30 == _myNewVec_35_T_3[5:0] ? myVec_48 : _GEN_1945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1947 = 6'h31 == _myNewVec_35_T_3[5:0] ? myVec_49 : _GEN_1946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1948 = 6'h32 == _myNewVec_35_T_3[5:0] ? myVec_50 : _GEN_1947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1949 = 6'h33 == _myNewVec_35_T_3[5:0] ? myVec_51 : _GEN_1948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1950 = 6'h34 == _myNewVec_35_T_3[5:0] ? myVec_52 : _GEN_1949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1951 = 6'h35 == _myNewVec_35_T_3[5:0] ? myVec_53 : _GEN_1950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1952 = 6'h36 == _myNewVec_35_T_3[5:0] ? myVec_54 : _GEN_1951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1953 = 6'h37 == _myNewVec_35_T_3[5:0] ? myVec_55 : _GEN_1952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1954 = 6'h38 == _myNewVec_35_T_3[5:0] ? myVec_56 : _GEN_1953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1955 = 6'h39 == _myNewVec_35_T_3[5:0] ? myVec_57 : _GEN_1954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1956 = 6'h3a == _myNewVec_35_T_3[5:0] ? myVec_58 : _GEN_1955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1957 = 6'h3b == _myNewVec_35_T_3[5:0] ? myVec_59 : _GEN_1956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1958 = 6'h3c == _myNewVec_35_T_3[5:0] ? myVec_60 : _GEN_1957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1959 = 6'h3d == _myNewVec_35_T_3[5:0] ? myVec_61 : _GEN_1958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1960 = 6'h3e == _myNewVec_35_T_3[5:0] ? myVec_62 : _GEN_1959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_35 = 6'h3f == _myNewVec_35_T_3[5:0] ? myVec_63 : _GEN_1960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_34_T_3 = _myNewVec_63_T_1 + 16'h1d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_1963 = 6'h1 == _myNewVec_34_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1964 = 6'h2 == _myNewVec_34_T_3[5:0] ? myVec_2 : _GEN_1963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1965 = 6'h3 == _myNewVec_34_T_3[5:0] ? myVec_3 : _GEN_1964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1966 = 6'h4 == _myNewVec_34_T_3[5:0] ? myVec_4 : _GEN_1965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1967 = 6'h5 == _myNewVec_34_T_3[5:0] ? myVec_5 : _GEN_1966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1968 = 6'h6 == _myNewVec_34_T_3[5:0] ? myVec_6 : _GEN_1967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1969 = 6'h7 == _myNewVec_34_T_3[5:0] ? myVec_7 : _GEN_1968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1970 = 6'h8 == _myNewVec_34_T_3[5:0] ? myVec_8 : _GEN_1969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1971 = 6'h9 == _myNewVec_34_T_3[5:0] ? myVec_9 : _GEN_1970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1972 = 6'ha == _myNewVec_34_T_3[5:0] ? myVec_10 : _GEN_1971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1973 = 6'hb == _myNewVec_34_T_3[5:0] ? myVec_11 : _GEN_1972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1974 = 6'hc == _myNewVec_34_T_3[5:0] ? myVec_12 : _GEN_1973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1975 = 6'hd == _myNewVec_34_T_3[5:0] ? myVec_13 : _GEN_1974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1976 = 6'he == _myNewVec_34_T_3[5:0] ? myVec_14 : _GEN_1975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1977 = 6'hf == _myNewVec_34_T_3[5:0] ? myVec_15 : _GEN_1976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1978 = 6'h10 == _myNewVec_34_T_3[5:0] ? myVec_16 : _GEN_1977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1979 = 6'h11 == _myNewVec_34_T_3[5:0] ? myVec_17 : _GEN_1978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1980 = 6'h12 == _myNewVec_34_T_3[5:0] ? myVec_18 : _GEN_1979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1981 = 6'h13 == _myNewVec_34_T_3[5:0] ? myVec_19 : _GEN_1980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1982 = 6'h14 == _myNewVec_34_T_3[5:0] ? myVec_20 : _GEN_1981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1983 = 6'h15 == _myNewVec_34_T_3[5:0] ? myVec_21 : _GEN_1982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1984 = 6'h16 == _myNewVec_34_T_3[5:0] ? myVec_22 : _GEN_1983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1985 = 6'h17 == _myNewVec_34_T_3[5:0] ? myVec_23 : _GEN_1984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1986 = 6'h18 == _myNewVec_34_T_3[5:0] ? myVec_24 : _GEN_1985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1987 = 6'h19 == _myNewVec_34_T_3[5:0] ? myVec_25 : _GEN_1986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1988 = 6'h1a == _myNewVec_34_T_3[5:0] ? myVec_26 : _GEN_1987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1989 = 6'h1b == _myNewVec_34_T_3[5:0] ? myVec_27 : _GEN_1988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1990 = 6'h1c == _myNewVec_34_T_3[5:0] ? myVec_28 : _GEN_1989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1991 = 6'h1d == _myNewVec_34_T_3[5:0] ? myVec_29 : _GEN_1990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1992 = 6'h1e == _myNewVec_34_T_3[5:0] ? myVec_30 : _GEN_1991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1993 = 6'h1f == _myNewVec_34_T_3[5:0] ? myVec_31 : _GEN_1992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1994 = 6'h20 == _myNewVec_34_T_3[5:0] ? myVec_32 : _GEN_1993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1995 = 6'h21 == _myNewVec_34_T_3[5:0] ? myVec_33 : _GEN_1994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1996 = 6'h22 == _myNewVec_34_T_3[5:0] ? myVec_34 : _GEN_1995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1997 = 6'h23 == _myNewVec_34_T_3[5:0] ? myVec_35 : _GEN_1996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1998 = 6'h24 == _myNewVec_34_T_3[5:0] ? myVec_36 : _GEN_1997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_1999 = 6'h25 == _myNewVec_34_T_3[5:0] ? myVec_37 : _GEN_1998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2000 = 6'h26 == _myNewVec_34_T_3[5:0] ? myVec_38 : _GEN_1999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2001 = 6'h27 == _myNewVec_34_T_3[5:0] ? myVec_39 : _GEN_2000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2002 = 6'h28 == _myNewVec_34_T_3[5:0] ? myVec_40 : _GEN_2001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2003 = 6'h29 == _myNewVec_34_T_3[5:0] ? myVec_41 : _GEN_2002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2004 = 6'h2a == _myNewVec_34_T_3[5:0] ? myVec_42 : _GEN_2003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2005 = 6'h2b == _myNewVec_34_T_3[5:0] ? myVec_43 : _GEN_2004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2006 = 6'h2c == _myNewVec_34_T_3[5:0] ? myVec_44 : _GEN_2005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2007 = 6'h2d == _myNewVec_34_T_3[5:0] ? myVec_45 : _GEN_2006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2008 = 6'h2e == _myNewVec_34_T_3[5:0] ? myVec_46 : _GEN_2007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2009 = 6'h2f == _myNewVec_34_T_3[5:0] ? myVec_47 : _GEN_2008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2010 = 6'h30 == _myNewVec_34_T_3[5:0] ? myVec_48 : _GEN_2009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2011 = 6'h31 == _myNewVec_34_T_3[5:0] ? myVec_49 : _GEN_2010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2012 = 6'h32 == _myNewVec_34_T_3[5:0] ? myVec_50 : _GEN_2011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2013 = 6'h33 == _myNewVec_34_T_3[5:0] ? myVec_51 : _GEN_2012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2014 = 6'h34 == _myNewVec_34_T_3[5:0] ? myVec_52 : _GEN_2013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2015 = 6'h35 == _myNewVec_34_T_3[5:0] ? myVec_53 : _GEN_2014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2016 = 6'h36 == _myNewVec_34_T_3[5:0] ? myVec_54 : _GEN_2015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2017 = 6'h37 == _myNewVec_34_T_3[5:0] ? myVec_55 : _GEN_2016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2018 = 6'h38 == _myNewVec_34_T_3[5:0] ? myVec_56 : _GEN_2017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2019 = 6'h39 == _myNewVec_34_T_3[5:0] ? myVec_57 : _GEN_2018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2020 = 6'h3a == _myNewVec_34_T_3[5:0] ? myVec_58 : _GEN_2019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2021 = 6'h3b == _myNewVec_34_T_3[5:0] ? myVec_59 : _GEN_2020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2022 = 6'h3c == _myNewVec_34_T_3[5:0] ? myVec_60 : _GEN_2021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2023 = 6'h3d == _myNewVec_34_T_3[5:0] ? myVec_61 : _GEN_2022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2024 = 6'h3e == _myNewVec_34_T_3[5:0] ? myVec_62 : _GEN_2023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_34 = 6'h3f == _myNewVec_34_T_3[5:0] ? myVec_63 : _GEN_2024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_33_T_3 = _myNewVec_63_T_1 + 16'h1e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2027 = 6'h1 == _myNewVec_33_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2028 = 6'h2 == _myNewVec_33_T_3[5:0] ? myVec_2 : _GEN_2027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2029 = 6'h3 == _myNewVec_33_T_3[5:0] ? myVec_3 : _GEN_2028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2030 = 6'h4 == _myNewVec_33_T_3[5:0] ? myVec_4 : _GEN_2029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2031 = 6'h5 == _myNewVec_33_T_3[5:0] ? myVec_5 : _GEN_2030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2032 = 6'h6 == _myNewVec_33_T_3[5:0] ? myVec_6 : _GEN_2031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2033 = 6'h7 == _myNewVec_33_T_3[5:0] ? myVec_7 : _GEN_2032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2034 = 6'h8 == _myNewVec_33_T_3[5:0] ? myVec_8 : _GEN_2033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2035 = 6'h9 == _myNewVec_33_T_3[5:0] ? myVec_9 : _GEN_2034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2036 = 6'ha == _myNewVec_33_T_3[5:0] ? myVec_10 : _GEN_2035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2037 = 6'hb == _myNewVec_33_T_3[5:0] ? myVec_11 : _GEN_2036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2038 = 6'hc == _myNewVec_33_T_3[5:0] ? myVec_12 : _GEN_2037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2039 = 6'hd == _myNewVec_33_T_3[5:0] ? myVec_13 : _GEN_2038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2040 = 6'he == _myNewVec_33_T_3[5:0] ? myVec_14 : _GEN_2039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2041 = 6'hf == _myNewVec_33_T_3[5:0] ? myVec_15 : _GEN_2040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2042 = 6'h10 == _myNewVec_33_T_3[5:0] ? myVec_16 : _GEN_2041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2043 = 6'h11 == _myNewVec_33_T_3[5:0] ? myVec_17 : _GEN_2042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2044 = 6'h12 == _myNewVec_33_T_3[5:0] ? myVec_18 : _GEN_2043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2045 = 6'h13 == _myNewVec_33_T_3[5:0] ? myVec_19 : _GEN_2044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2046 = 6'h14 == _myNewVec_33_T_3[5:0] ? myVec_20 : _GEN_2045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2047 = 6'h15 == _myNewVec_33_T_3[5:0] ? myVec_21 : _GEN_2046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2048 = 6'h16 == _myNewVec_33_T_3[5:0] ? myVec_22 : _GEN_2047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2049 = 6'h17 == _myNewVec_33_T_3[5:0] ? myVec_23 : _GEN_2048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2050 = 6'h18 == _myNewVec_33_T_3[5:0] ? myVec_24 : _GEN_2049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2051 = 6'h19 == _myNewVec_33_T_3[5:0] ? myVec_25 : _GEN_2050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2052 = 6'h1a == _myNewVec_33_T_3[5:0] ? myVec_26 : _GEN_2051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2053 = 6'h1b == _myNewVec_33_T_3[5:0] ? myVec_27 : _GEN_2052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2054 = 6'h1c == _myNewVec_33_T_3[5:0] ? myVec_28 : _GEN_2053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2055 = 6'h1d == _myNewVec_33_T_3[5:0] ? myVec_29 : _GEN_2054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2056 = 6'h1e == _myNewVec_33_T_3[5:0] ? myVec_30 : _GEN_2055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2057 = 6'h1f == _myNewVec_33_T_3[5:0] ? myVec_31 : _GEN_2056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2058 = 6'h20 == _myNewVec_33_T_3[5:0] ? myVec_32 : _GEN_2057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2059 = 6'h21 == _myNewVec_33_T_3[5:0] ? myVec_33 : _GEN_2058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2060 = 6'h22 == _myNewVec_33_T_3[5:0] ? myVec_34 : _GEN_2059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2061 = 6'h23 == _myNewVec_33_T_3[5:0] ? myVec_35 : _GEN_2060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2062 = 6'h24 == _myNewVec_33_T_3[5:0] ? myVec_36 : _GEN_2061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2063 = 6'h25 == _myNewVec_33_T_3[5:0] ? myVec_37 : _GEN_2062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2064 = 6'h26 == _myNewVec_33_T_3[5:0] ? myVec_38 : _GEN_2063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2065 = 6'h27 == _myNewVec_33_T_3[5:0] ? myVec_39 : _GEN_2064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2066 = 6'h28 == _myNewVec_33_T_3[5:0] ? myVec_40 : _GEN_2065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2067 = 6'h29 == _myNewVec_33_T_3[5:0] ? myVec_41 : _GEN_2066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2068 = 6'h2a == _myNewVec_33_T_3[5:0] ? myVec_42 : _GEN_2067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2069 = 6'h2b == _myNewVec_33_T_3[5:0] ? myVec_43 : _GEN_2068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2070 = 6'h2c == _myNewVec_33_T_3[5:0] ? myVec_44 : _GEN_2069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2071 = 6'h2d == _myNewVec_33_T_3[5:0] ? myVec_45 : _GEN_2070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2072 = 6'h2e == _myNewVec_33_T_3[5:0] ? myVec_46 : _GEN_2071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2073 = 6'h2f == _myNewVec_33_T_3[5:0] ? myVec_47 : _GEN_2072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2074 = 6'h30 == _myNewVec_33_T_3[5:0] ? myVec_48 : _GEN_2073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2075 = 6'h31 == _myNewVec_33_T_3[5:0] ? myVec_49 : _GEN_2074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2076 = 6'h32 == _myNewVec_33_T_3[5:0] ? myVec_50 : _GEN_2075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2077 = 6'h33 == _myNewVec_33_T_3[5:0] ? myVec_51 : _GEN_2076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2078 = 6'h34 == _myNewVec_33_T_3[5:0] ? myVec_52 : _GEN_2077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2079 = 6'h35 == _myNewVec_33_T_3[5:0] ? myVec_53 : _GEN_2078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2080 = 6'h36 == _myNewVec_33_T_3[5:0] ? myVec_54 : _GEN_2079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2081 = 6'h37 == _myNewVec_33_T_3[5:0] ? myVec_55 : _GEN_2080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2082 = 6'h38 == _myNewVec_33_T_3[5:0] ? myVec_56 : _GEN_2081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2083 = 6'h39 == _myNewVec_33_T_3[5:0] ? myVec_57 : _GEN_2082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2084 = 6'h3a == _myNewVec_33_T_3[5:0] ? myVec_58 : _GEN_2083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2085 = 6'h3b == _myNewVec_33_T_3[5:0] ? myVec_59 : _GEN_2084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2086 = 6'h3c == _myNewVec_33_T_3[5:0] ? myVec_60 : _GEN_2085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2087 = 6'h3d == _myNewVec_33_T_3[5:0] ? myVec_61 : _GEN_2086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2088 = 6'h3e == _myNewVec_33_T_3[5:0] ? myVec_62 : _GEN_2087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_33 = 6'h3f == _myNewVec_33_T_3[5:0] ? myVec_63 : _GEN_2088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_32_T_3 = _myNewVec_63_T_1 + 16'h1f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2091 = 6'h1 == _myNewVec_32_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2092 = 6'h2 == _myNewVec_32_T_3[5:0] ? myVec_2 : _GEN_2091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2093 = 6'h3 == _myNewVec_32_T_3[5:0] ? myVec_3 : _GEN_2092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2094 = 6'h4 == _myNewVec_32_T_3[5:0] ? myVec_4 : _GEN_2093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2095 = 6'h5 == _myNewVec_32_T_3[5:0] ? myVec_5 : _GEN_2094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2096 = 6'h6 == _myNewVec_32_T_3[5:0] ? myVec_6 : _GEN_2095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2097 = 6'h7 == _myNewVec_32_T_3[5:0] ? myVec_7 : _GEN_2096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2098 = 6'h8 == _myNewVec_32_T_3[5:0] ? myVec_8 : _GEN_2097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2099 = 6'h9 == _myNewVec_32_T_3[5:0] ? myVec_9 : _GEN_2098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2100 = 6'ha == _myNewVec_32_T_3[5:0] ? myVec_10 : _GEN_2099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2101 = 6'hb == _myNewVec_32_T_3[5:0] ? myVec_11 : _GEN_2100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2102 = 6'hc == _myNewVec_32_T_3[5:0] ? myVec_12 : _GEN_2101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2103 = 6'hd == _myNewVec_32_T_3[5:0] ? myVec_13 : _GEN_2102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2104 = 6'he == _myNewVec_32_T_3[5:0] ? myVec_14 : _GEN_2103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2105 = 6'hf == _myNewVec_32_T_3[5:0] ? myVec_15 : _GEN_2104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2106 = 6'h10 == _myNewVec_32_T_3[5:0] ? myVec_16 : _GEN_2105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2107 = 6'h11 == _myNewVec_32_T_3[5:0] ? myVec_17 : _GEN_2106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2108 = 6'h12 == _myNewVec_32_T_3[5:0] ? myVec_18 : _GEN_2107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2109 = 6'h13 == _myNewVec_32_T_3[5:0] ? myVec_19 : _GEN_2108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2110 = 6'h14 == _myNewVec_32_T_3[5:0] ? myVec_20 : _GEN_2109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2111 = 6'h15 == _myNewVec_32_T_3[5:0] ? myVec_21 : _GEN_2110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2112 = 6'h16 == _myNewVec_32_T_3[5:0] ? myVec_22 : _GEN_2111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2113 = 6'h17 == _myNewVec_32_T_3[5:0] ? myVec_23 : _GEN_2112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2114 = 6'h18 == _myNewVec_32_T_3[5:0] ? myVec_24 : _GEN_2113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2115 = 6'h19 == _myNewVec_32_T_3[5:0] ? myVec_25 : _GEN_2114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2116 = 6'h1a == _myNewVec_32_T_3[5:0] ? myVec_26 : _GEN_2115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2117 = 6'h1b == _myNewVec_32_T_3[5:0] ? myVec_27 : _GEN_2116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2118 = 6'h1c == _myNewVec_32_T_3[5:0] ? myVec_28 : _GEN_2117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2119 = 6'h1d == _myNewVec_32_T_3[5:0] ? myVec_29 : _GEN_2118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2120 = 6'h1e == _myNewVec_32_T_3[5:0] ? myVec_30 : _GEN_2119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2121 = 6'h1f == _myNewVec_32_T_3[5:0] ? myVec_31 : _GEN_2120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2122 = 6'h20 == _myNewVec_32_T_3[5:0] ? myVec_32 : _GEN_2121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2123 = 6'h21 == _myNewVec_32_T_3[5:0] ? myVec_33 : _GEN_2122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2124 = 6'h22 == _myNewVec_32_T_3[5:0] ? myVec_34 : _GEN_2123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2125 = 6'h23 == _myNewVec_32_T_3[5:0] ? myVec_35 : _GEN_2124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2126 = 6'h24 == _myNewVec_32_T_3[5:0] ? myVec_36 : _GEN_2125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2127 = 6'h25 == _myNewVec_32_T_3[5:0] ? myVec_37 : _GEN_2126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2128 = 6'h26 == _myNewVec_32_T_3[5:0] ? myVec_38 : _GEN_2127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2129 = 6'h27 == _myNewVec_32_T_3[5:0] ? myVec_39 : _GEN_2128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2130 = 6'h28 == _myNewVec_32_T_3[5:0] ? myVec_40 : _GEN_2129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2131 = 6'h29 == _myNewVec_32_T_3[5:0] ? myVec_41 : _GEN_2130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2132 = 6'h2a == _myNewVec_32_T_3[5:0] ? myVec_42 : _GEN_2131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2133 = 6'h2b == _myNewVec_32_T_3[5:0] ? myVec_43 : _GEN_2132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2134 = 6'h2c == _myNewVec_32_T_3[5:0] ? myVec_44 : _GEN_2133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2135 = 6'h2d == _myNewVec_32_T_3[5:0] ? myVec_45 : _GEN_2134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2136 = 6'h2e == _myNewVec_32_T_3[5:0] ? myVec_46 : _GEN_2135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2137 = 6'h2f == _myNewVec_32_T_3[5:0] ? myVec_47 : _GEN_2136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2138 = 6'h30 == _myNewVec_32_T_3[5:0] ? myVec_48 : _GEN_2137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2139 = 6'h31 == _myNewVec_32_T_3[5:0] ? myVec_49 : _GEN_2138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2140 = 6'h32 == _myNewVec_32_T_3[5:0] ? myVec_50 : _GEN_2139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2141 = 6'h33 == _myNewVec_32_T_3[5:0] ? myVec_51 : _GEN_2140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2142 = 6'h34 == _myNewVec_32_T_3[5:0] ? myVec_52 : _GEN_2141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2143 = 6'h35 == _myNewVec_32_T_3[5:0] ? myVec_53 : _GEN_2142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2144 = 6'h36 == _myNewVec_32_T_3[5:0] ? myVec_54 : _GEN_2143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2145 = 6'h37 == _myNewVec_32_T_3[5:0] ? myVec_55 : _GEN_2144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2146 = 6'h38 == _myNewVec_32_T_3[5:0] ? myVec_56 : _GEN_2145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2147 = 6'h39 == _myNewVec_32_T_3[5:0] ? myVec_57 : _GEN_2146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2148 = 6'h3a == _myNewVec_32_T_3[5:0] ? myVec_58 : _GEN_2147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2149 = 6'h3b == _myNewVec_32_T_3[5:0] ? myVec_59 : _GEN_2148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2150 = 6'h3c == _myNewVec_32_T_3[5:0] ? myVec_60 : _GEN_2149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2151 = 6'h3d == _myNewVec_32_T_3[5:0] ? myVec_61 : _GEN_2150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2152 = 6'h3e == _myNewVec_32_T_3[5:0] ? myVec_62 : _GEN_2151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_32 = 6'h3f == _myNewVec_32_T_3[5:0] ? myVec_63 : _GEN_2152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_hi_lo_lo = {myNewVec_39,myNewVec_38,myNewVec_37,myNewVec_36,myNewVec_35,myNewVec_34,myNewVec_33
    ,myNewVec_32}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_hi_lo = {myNewVec_47,myNewVec_46,myNewVec_45,myNewVec_44,myNewVec_43,myNewVec_42,myNewVec_41,
    myNewVec_40,myNewWire_hi_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_hi = {myNewVec_63,myNewVec_62,myNewVec_61,myNewVec_60,myNewVec_59,myNewVec_58,myNewVec_57,
    myNewVec_56,myNewWire_hi_hi_lo,myNewWire_hi_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_31_T_3 = _myNewVec_63_T_1 + 16'h20; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2155 = 6'h1 == _myNewVec_31_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2156 = 6'h2 == _myNewVec_31_T_3[5:0] ? myVec_2 : _GEN_2155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2157 = 6'h3 == _myNewVec_31_T_3[5:0] ? myVec_3 : _GEN_2156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2158 = 6'h4 == _myNewVec_31_T_3[5:0] ? myVec_4 : _GEN_2157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2159 = 6'h5 == _myNewVec_31_T_3[5:0] ? myVec_5 : _GEN_2158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2160 = 6'h6 == _myNewVec_31_T_3[5:0] ? myVec_6 : _GEN_2159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2161 = 6'h7 == _myNewVec_31_T_3[5:0] ? myVec_7 : _GEN_2160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2162 = 6'h8 == _myNewVec_31_T_3[5:0] ? myVec_8 : _GEN_2161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2163 = 6'h9 == _myNewVec_31_T_3[5:0] ? myVec_9 : _GEN_2162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2164 = 6'ha == _myNewVec_31_T_3[5:0] ? myVec_10 : _GEN_2163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2165 = 6'hb == _myNewVec_31_T_3[5:0] ? myVec_11 : _GEN_2164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2166 = 6'hc == _myNewVec_31_T_3[5:0] ? myVec_12 : _GEN_2165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2167 = 6'hd == _myNewVec_31_T_3[5:0] ? myVec_13 : _GEN_2166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2168 = 6'he == _myNewVec_31_T_3[5:0] ? myVec_14 : _GEN_2167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2169 = 6'hf == _myNewVec_31_T_3[5:0] ? myVec_15 : _GEN_2168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2170 = 6'h10 == _myNewVec_31_T_3[5:0] ? myVec_16 : _GEN_2169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2171 = 6'h11 == _myNewVec_31_T_3[5:0] ? myVec_17 : _GEN_2170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2172 = 6'h12 == _myNewVec_31_T_3[5:0] ? myVec_18 : _GEN_2171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2173 = 6'h13 == _myNewVec_31_T_3[5:0] ? myVec_19 : _GEN_2172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2174 = 6'h14 == _myNewVec_31_T_3[5:0] ? myVec_20 : _GEN_2173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2175 = 6'h15 == _myNewVec_31_T_3[5:0] ? myVec_21 : _GEN_2174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2176 = 6'h16 == _myNewVec_31_T_3[5:0] ? myVec_22 : _GEN_2175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2177 = 6'h17 == _myNewVec_31_T_3[5:0] ? myVec_23 : _GEN_2176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2178 = 6'h18 == _myNewVec_31_T_3[5:0] ? myVec_24 : _GEN_2177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2179 = 6'h19 == _myNewVec_31_T_3[5:0] ? myVec_25 : _GEN_2178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2180 = 6'h1a == _myNewVec_31_T_3[5:0] ? myVec_26 : _GEN_2179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2181 = 6'h1b == _myNewVec_31_T_3[5:0] ? myVec_27 : _GEN_2180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2182 = 6'h1c == _myNewVec_31_T_3[5:0] ? myVec_28 : _GEN_2181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2183 = 6'h1d == _myNewVec_31_T_3[5:0] ? myVec_29 : _GEN_2182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2184 = 6'h1e == _myNewVec_31_T_3[5:0] ? myVec_30 : _GEN_2183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2185 = 6'h1f == _myNewVec_31_T_3[5:0] ? myVec_31 : _GEN_2184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2186 = 6'h20 == _myNewVec_31_T_3[5:0] ? myVec_32 : _GEN_2185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2187 = 6'h21 == _myNewVec_31_T_3[5:0] ? myVec_33 : _GEN_2186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2188 = 6'h22 == _myNewVec_31_T_3[5:0] ? myVec_34 : _GEN_2187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2189 = 6'h23 == _myNewVec_31_T_3[5:0] ? myVec_35 : _GEN_2188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2190 = 6'h24 == _myNewVec_31_T_3[5:0] ? myVec_36 : _GEN_2189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2191 = 6'h25 == _myNewVec_31_T_3[5:0] ? myVec_37 : _GEN_2190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2192 = 6'h26 == _myNewVec_31_T_3[5:0] ? myVec_38 : _GEN_2191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2193 = 6'h27 == _myNewVec_31_T_3[5:0] ? myVec_39 : _GEN_2192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2194 = 6'h28 == _myNewVec_31_T_3[5:0] ? myVec_40 : _GEN_2193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2195 = 6'h29 == _myNewVec_31_T_3[5:0] ? myVec_41 : _GEN_2194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2196 = 6'h2a == _myNewVec_31_T_3[5:0] ? myVec_42 : _GEN_2195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2197 = 6'h2b == _myNewVec_31_T_3[5:0] ? myVec_43 : _GEN_2196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2198 = 6'h2c == _myNewVec_31_T_3[5:0] ? myVec_44 : _GEN_2197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2199 = 6'h2d == _myNewVec_31_T_3[5:0] ? myVec_45 : _GEN_2198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2200 = 6'h2e == _myNewVec_31_T_3[5:0] ? myVec_46 : _GEN_2199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2201 = 6'h2f == _myNewVec_31_T_3[5:0] ? myVec_47 : _GEN_2200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2202 = 6'h30 == _myNewVec_31_T_3[5:0] ? myVec_48 : _GEN_2201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2203 = 6'h31 == _myNewVec_31_T_3[5:0] ? myVec_49 : _GEN_2202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2204 = 6'h32 == _myNewVec_31_T_3[5:0] ? myVec_50 : _GEN_2203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2205 = 6'h33 == _myNewVec_31_T_3[5:0] ? myVec_51 : _GEN_2204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2206 = 6'h34 == _myNewVec_31_T_3[5:0] ? myVec_52 : _GEN_2205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2207 = 6'h35 == _myNewVec_31_T_3[5:0] ? myVec_53 : _GEN_2206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2208 = 6'h36 == _myNewVec_31_T_3[5:0] ? myVec_54 : _GEN_2207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2209 = 6'h37 == _myNewVec_31_T_3[5:0] ? myVec_55 : _GEN_2208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2210 = 6'h38 == _myNewVec_31_T_3[5:0] ? myVec_56 : _GEN_2209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2211 = 6'h39 == _myNewVec_31_T_3[5:0] ? myVec_57 : _GEN_2210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2212 = 6'h3a == _myNewVec_31_T_3[5:0] ? myVec_58 : _GEN_2211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2213 = 6'h3b == _myNewVec_31_T_3[5:0] ? myVec_59 : _GEN_2212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2214 = 6'h3c == _myNewVec_31_T_3[5:0] ? myVec_60 : _GEN_2213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2215 = 6'h3d == _myNewVec_31_T_3[5:0] ? myVec_61 : _GEN_2214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2216 = 6'h3e == _myNewVec_31_T_3[5:0] ? myVec_62 : _GEN_2215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_31 = 6'h3f == _myNewVec_31_T_3[5:0] ? myVec_63 : _GEN_2216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_30_T_3 = _myNewVec_63_T_1 + 16'h21; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2219 = 6'h1 == _myNewVec_30_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2220 = 6'h2 == _myNewVec_30_T_3[5:0] ? myVec_2 : _GEN_2219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2221 = 6'h3 == _myNewVec_30_T_3[5:0] ? myVec_3 : _GEN_2220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2222 = 6'h4 == _myNewVec_30_T_3[5:0] ? myVec_4 : _GEN_2221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2223 = 6'h5 == _myNewVec_30_T_3[5:0] ? myVec_5 : _GEN_2222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2224 = 6'h6 == _myNewVec_30_T_3[5:0] ? myVec_6 : _GEN_2223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2225 = 6'h7 == _myNewVec_30_T_3[5:0] ? myVec_7 : _GEN_2224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2226 = 6'h8 == _myNewVec_30_T_3[5:0] ? myVec_8 : _GEN_2225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2227 = 6'h9 == _myNewVec_30_T_3[5:0] ? myVec_9 : _GEN_2226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2228 = 6'ha == _myNewVec_30_T_3[5:0] ? myVec_10 : _GEN_2227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2229 = 6'hb == _myNewVec_30_T_3[5:0] ? myVec_11 : _GEN_2228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2230 = 6'hc == _myNewVec_30_T_3[5:0] ? myVec_12 : _GEN_2229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2231 = 6'hd == _myNewVec_30_T_3[5:0] ? myVec_13 : _GEN_2230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2232 = 6'he == _myNewVec_30_T_3[5:0] ? myVec_14 : _GEN_2231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2233 = 6'hf == _myNewVec_30_T_3[5:0] ? myVec_15 : _GEN_2232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2234 = 6'h10 == _myNewVec_30_T_3[5:0] ? myVec_16 : _GEN_2233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2235 = 6'h11 == _myNewVec_30_T_3[5:0] ? myVec_17 : _GEN_2234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2236 = 6'h12 == _myNewVec_30_T_3[5:0] ? myVec_18 : _GEN_2235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2237 = 6'h13 == _myNewVec_30_T_3[5:0] ? myVec_19 : _GEN_2236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2238 = 6'h14 == _myNewVec_30_T_3[5:0] ? myVec_20 : _GEN_2237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2239 = 6'h15 == _myNewVec_30_T_3[5:0] ? myVec_21 : _GEN_2238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2240 = 6'h16 == _myNewVec_30_T_3[5:0] ? myVec_22 : _GEN_2239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2241 = 6'h17 == _myNewVec_30_T_3[5:0] ? myVec_23 : _GEN_2240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2242 = 6'h18 == _myNewVec_30_T_3[5:0] ? myVec_24 : _GEN_2241; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2243 = 6'h19 == _myNewVec_30_T_3[5:0] ? myVec_25 : _GEN_2242; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2244 = 6'h1a == _myNewVec_30_T_3[5:0] ? myVec_26 : _GEN_2243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2245 = 6'h1b == _myNewVec_30_T_3[5:0] ? myVec_27 : _GEN_2244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2246 = 6'h1c == _myNewVec_30_T_3[5:0] ? myVec_28 : _GEN_2245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2247 = 6'h1d == _myNewVec_30_T_3[5:0] ? myVec_29 : _GEN_2246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2248 = 6'h1e == _myNewVec_30_T_3[5:0] ? myVec_30 : _GEN_2247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2249 = 6'h1f == _myNewVec_30_T_3[5:0] ? myVec_31 : _GEN_2248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2250 = 6'h20 == _myNewVec_30_T_3[5:0] ? myVec_32 : _GEN_2249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2251 = 6'h21 == _myNewVec_30_T_3[5:0] ? myVec_33 : _GEN_2250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2252 = 6'h22 == _myNewVec_30_T_3[5:0] ? myVec_34 : _GEN_2251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2253 = 6'h23 == _myNewVec_30_T_3[5:0] ? myVec_35 : _GEN_2252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2254 = 6'h24 == _myNewVec_30_T_3[5:0] ? myVec_36 : _GEN_2253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2255 = 6'h25 == _myNewVec_30_T_3[5:0] ? myVec_37 : _GEN_2254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2256 = 6'h26 == _myNewVec_30_T_3[5:0] ? myVec_38 : _GEN_2255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2257 = 6'h27 == _myNewVec_30_T_3[5:0] ? myVec_39 : _GEN_2256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2258 = 6'h28 == _myNewVec_30_T_3[5:0] ? myVec_40 : _GEN_2257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2259 = 6'h29 == _myNewVec_30_T_3[5:0] ? myVec_41 : _GEN_2258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2260 = 6'h2a == _myNewVec_30_T_3[5:0] ? myVec_42 : _GEN_2259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2261 = 6'h2b == _myNewVec_30_T_3[5:0] ? myVec_43 : _GEN_2260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2262 = 6'h2c == _myNewVec_30_T_3[5:0] ? myVec_44 : _GEN_2261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2263 = 6'h2d == _myNewVec_30_T_3[5:0] ? myVec_45 : _GEN_2262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2264 = 6'h2e == _myNewVec_30_T_3[5:0] ? myVec_46 : _GEN_2263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2265 = 6'h2f == _myNewVec_30_T_3[5:0] ? myVec_47 : _GEN_2264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2266 = 6'h30 == _myNewVec_30_T_3[5:0] ? myVec_48 : _GEN_2265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2267 = 6'h31 == _myNewVec_30_T_3[5:0] ? myVec_49 : _GEN_2266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2268 = 6'h32 == _myNewVec_30_T_3[5:0] ? myVec_50 : _GEN_2267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2269 = 6'h33 == _myNewVec_30_T_3[5:0] ? myVec_51 : _GEN_2268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2270 = 6'h34 == _myNewVec_30_T_3[5:0] ? myVec_52 : _GEN_2269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2271 = 6'h35 == _myNewVec_30_T_3[5:0] ? myVec_53 : _GEN_2270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2272 = 6'h36 == _myNewVec_30_T_3[5:0] ? myVec_54 : _GEN_2271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2273 = 6'h37 == _myNewVec_30_T_3[5:0] ? myVec_55 : _GEN_2272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2274 = 6'h38 == _myNewVec_30_T_3[5:0] ? myVec_56 : _GEN_2273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2275 = 6'h39 == _myNewVec_30_T_3[5:0] ? myVec_57 : _GEN_2274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2276 = 6'h3a == _myNewVec_30_T_3[5:0] ? myVec_58 : _GEN_2275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2277 = 6'h3b == _myNewVec_30_T_3[5:0] ? myVec_59 : _GEN_2276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2278 = 6'h3c == _myNewVec_30_T_3[5:0] ? myVec_60 : _GEN_2277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2279 = 6'h3d == _myNewVec_30_T_3[5:0] ? myVec_61 : _GEN_2278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2280 = 6'h3e == _myNewVec_30_T_3[5:0] ? myVec_62 : _GEN_2279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_30 = 6'h3f == _myNewVec_30_T_3[5:0] ? myVec_63 : _GEN_2280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_29_T_3 = _myNewVec_63_T_1 + 16'h22; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2283 = 6'h1 == _myNewVec_29_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2284 = 6'h2 == _myNewVec_29_T_3[5:0] ? myVec_2 : _GEN_2283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2285 = 6'h3 == _myNewVec_29_T_3[5:0] ? myVec_3 : _GEN_2284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2286 = 6'h4 == _myNewVec_29_T_3[5:0] ? myVec_4 : _GEN_2285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2287 = 6'h5 == _myNewVec_29_T_3[5:0] ? myVec_5 : _GEN_2286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2288 = 6'h6 == _myNewVec_29_T_3[5:0] ? myVec_6 : _GEN_2287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2289 = 6'h7 == _myNewVec_29_T_3[5:0] ? myVec_7 : _GEN_2288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2290 = 6'h8 == _myNewVec_29_T_3[5:0] ? myVec_8 : _GEN_2289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2291 = 6'h9 == _myNewVec_29_T_3[5:0] ? myVec_9 : _GEN_2290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2292 = 6'ha == _myNewVec_29_T_3[5:0] ? myVec_10 : _GEN_2291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2293 = 6'hb == _myNewVec_29_T_3[5:0] ? myVec_11 : _GEN_2292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2294 = 6'hc == _myNewVec_29_T_3[5:0] ? myVec_12 : _GEN_2293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2295 = 6'hd == _myNewVec_29_T_3[5:0] ? myVec_13 : _GEN_2294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2296 = 6'he == _myNewVec_29_T_3[5:0] ? myVec_14 : _GEN_2295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2297 = 6'hf == _myNewVec_29_T_3[5:0] ? myVec_15 : _GEN_2296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2298 = 6'h10 == _myNewVec_29_T_3[5:0] ? myVec_16 : _GEN_2297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2299 = 6'h11 == _myNewVec_29_T_3[5:0] ? myVec_17 : _GEN_2298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2300 = 6'h12 == _myNewVec_29_T_3[5:0] ? myVec_18 : _GEN_2299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2301 = 6'h13 == _myNewVec_29_T_3[5:0] ? myVec_19 : _GEN_2300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2302 = 6'h14 == _myNewVec_29_T_3[5:0] ? myVec_20 : _GEN_2301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2303 = 6'h15 == _myNewVec_29_T_3[5:0] ? myVec_21 : _GEN_2302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2304 = 6'h16 == _myNewVec_29_T_3[5:0] ? myVec_22 : _GEN_2303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2305 = 6'h17 == _myNewVec_29_T_3[5:0] ? myVec_23 : _GEN_2304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2306 = 6'h18 == _myNewVec_29_T_3[5:0] ? myVec_24 : _GEN_2305; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2307 = 6'h19 == _myNewVec_29_T_3[5:0] ? myVec_25 : _GEN_2306; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2308 = 6'h1a == _myNewVec_29_T_3[5:0] ? myVec_26 : _GEN_2307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2309 = 6'h1b == _myNewVec_29_T_3[5:0] ? myVec_27 : _GEN_2308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2310 = 6'h1c == _myNewVec_29_T_3[5:0] ? myVec_28 : _GEN_2309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2311 = 6'h1d == _myNewVec_29_T_3[5:0] ? myVec_29 : _GEN_2310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2312 = 6'h1e == _myNewVec_29_T_3[5:0] ? myVec_30 : _GEN_2311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2313 = 6'h1f == _myNewVec_29_T_3[5:0] ? myVec_31 : _GEN_2312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2314 = 6'h20 == _myNewVec_29_T_3[5:0] ? myVec_32 : _GEN_2313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2315 = 6'h21 == _myNewVec_29_T_3[5:0] ? myVec_33 : _GEN_2314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2316 = 6'h22 == _myNewVec_29_T_3[5:0] ? myVec_34 : _GEN_2315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2317 = 6'h23 == _myNewVec_29_T_3[5:0] ? myVec_35 : _GEN_2316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2318 = 6'h24 == _myNewVec_29_T_3[5:0] ? myVec_36 : _GEN_2317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2319 = 6'h25 == _myNewVec_29_T_3[5:0] ? myVec_37 : _GEN_2318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2320 = 6'h26 == _myNewVec_29_T_3[5:0] ? myVec_38 : _GEN_2319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2321 = 6'h27 == _myNewVec_29_T_3[5:0] ? myVec_39 : _GEN_2320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2322 = 6'h28 == _myNewVec_29_T_3[5:0] ? myVec_40 : _GEN_2321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2323 = 6'h29 == _myNewVec_29_T_3[5:0] ? myVec_41 : _GEN_2322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2324 = 6'h2a == _myNewVec_29_T_3[5:0] ? myVec_42 : _GEN_2323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2325 = 6'h2b == _myNewVec_29_T_3[5:0] ? myVec_43 : _GEN_2324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2326 = 6'h2c == _myNewVec_29_T_3[5:0] ? myVec_44 : _GEN_2325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2327 = 6'h2d == _myNewVec_29_T_3[5:0] ? myVec_45 : _GEN_2326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2328 = 6'h2e == _myNewVec_29_T_3[5:0] ? myVec_46 : _GEN_2327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2329 = 6'h2f == _myNewVec_29_T_3[5:0] ? myVec_47 : _GEN_2328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2330 = 6'h30 == _myNewVec_29_T_3[5:0] ? myVec_48 : _GEN_2329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2331 = 6'h31 == _myNewVec_29_T_3[5:0] ? myVec_49 : _GEN_2330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2332 = 6'h32 == _myNewVec_29_T_3[5:0] ? myVec_50 : _GEN_2331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2333 = 6'h33 == _myNewVec_29_T_3[5:0] ? myVec_51 : _GEN_2332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2334 = 6'h34 == _myNewVec_29_T_3[5:0] ? myVec_52 : _GEN_2333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2335 = 6'h35 == _myNewVec_29_T_3[5:0] ? myVec_53 : _GEN_2334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2336 = 6'h36 == _myNewVec_29_T_3[5:0] ? myVec_54 : _GEN_2335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2337 = 6'h37 == _myNewVec_29_T_3[5:0] ? myVec_55 : _GEN_2336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2338 = 6'h38 == _myNewVec_29_T_3[5:0] ? myVec_56 : _GEN_2337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2339 = 6'h39 == _myNewVec_29_T_3[5:0] ? myVec_57 : _GEN_2338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2340 = 6'h3a == _myNewVec_29_T_3[5:0] ? myVec_58 : _GEN_2339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2341 = 6'h3b == _myNewVec_29_T_3[5:0] ? myVec_59 : _GEN_2340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2342 = 6'h3c == _myNewVec_29_T_3[5:0] ? myVec_60 : _GEN_2341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2343 = 6'h3d == _myNewVec_29_T_3[5:0] ? myVec_61 : _GEN_2342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2344 = 6'h3e == _myNewVec_29_T_3[5:0] ? myVec_62 : _GEN_2343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_29 = 6'h3f == _myNewVec_29_T_3[5:0] ? myVec_63 : _GEN_2344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_28_T_3 = _myNewVec_63_T_1 + 16'h23; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2347 = 6'h1 == _myNewVec_28_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2348 = 6'h2 == _myNewVec_28_T_3[5:0] ? myVec_2 : _GEN_2347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2349 = 6'h3 == _myNewVec_28_T_3[5:0] ? myVec_3 : _GEN_2348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2350 = 6'h4 == _myNewVec_28_T_3[5:0] ? myVec_4 : _GEN_2349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2351 = 6'h5 == _myNewVec_28_T_3[5:0] ? myVec_5 : _GEN_2350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2352 = 6'h6 == _myNewVec_28_T_3[5:0] ? myVec_6 : _GEN_2351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2353 = 6'h7 == _myNewVec_28_T_3[5:0] ? myVec_7 : _GEN_2352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2354 = 6'h8 == _myNewVec_28_T_3[5:0] ? myVec_8 : _GEN_2353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2355 = 6'h9 == _myNewVec_28_T_3[5:0] ? myVec_9 : _GEN_2354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2356 = 6'ha == _myNewVec_28_T_3[5:0] ? myVec_10 : _GEN_2355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2357 = 6'hb == _myNewVec_28_T_3[5:0] ? myVec_11 : _GEN_2356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2358 = 6'hc == _myNewVec_28_T_3[5:0] ? myVec_12 : _GEN_2357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2359 = 6'hd == _myNewVec_28_T_3[5:0] ? myVec_13 : _GEN_2358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2360 = 6'he == _myNewVec_28_T_3[5:0] ? myVec_14 : _GEN_2359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2361 = 6'hf == _myNewVec_28_T_3[5:0] ? myVec_15 : _GEN_2360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2362 = 6'h10 == _myNewVec_28_T_3[5:0] ? myVec_16 : _GEN_2361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2363 = 6'h11 == _myNewVec_28_T_3[5:0] ? myVec_17 : _GEN_2362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2364 = 6'h12 == _myNewVec_28_T_3[5:0] ? myVec_18 : _GEN_2363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2365 = 6'h13 == _myNewVec_28_T_3[5:0] ? myVec_19 : _GEN_2364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2366 = 6'h14 == _myNewVec_28_T_3[5:0] ? myVec_20 : _GEN_2365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2367 = 6'h15 == _myNewVec_28_T_3[5:0] ? myVec_21 : _GEN_2366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2368 = 6'h16 == _myNewVec_28_T_3[5:0] ? myVec_22 : _GEN_2367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2369 = 6'h17 == _myNewVec_28_T_3[5:0] ? myVec_23 : _GEN_2368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2370 = 6'h18 == _myNewVec_28_T_3[5:0] ? myVec_24 : _GEN_2369; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2371 = 6'h19 == _myNewVec_28_T_3[5:0] ? myVec_25 : _GEN_2370; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2372 = 6'h1a == _myNewVec_28_T_3[5:0] ? myVec_26 : _GEN_2371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2373 = 6'h1b == _myNewVec_28_T_3[5:0] ? myVec_27 : _GEN_2372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2374 = 6'h1c == _myNewVec_28_T_3[5:0] ? myVec_28 : _GEN_2373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2375 = 6'h1d == _myNewVec_28_T_3[5:0] ? myVec_29 : _GEN_2374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2376 = 6'h1e == _myNewVec_28_T_3[5:0] ? myVec_30 : _GEN_2375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2377 = 6'h1f == _myNewVec_28_T_3[5:0] ? myVec_31 : _GEN_2376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2378 = 6'h20 == _myNewVec_28_T_3[5:0] ? myVec_32 : _GEN_2377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2379 = 6'h21 == _myNewVec_28_T_3[5:0] ? myVec_33 : _GEN_2378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2380 = 6'h22 == _myNewVec_28_T_3[5:0] ? myVec_34 : _GEN_2379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2381 = 6'h23 == _myNewVec_28_T_3[5:0] ? myVec_35 : _GEN_2380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2382 = 6'h24 == _myNewVec_28_T_3[5:0] ? myVec_36 : _GEN_2381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2383 = 6'h25 == _myNewVec_28_T_3[5:0] ? myVec_37 : _GEN_2382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2384 = 6'h26 == _myNewVec_28_T_3[5:0] ? myVec_38 : _GEN_2383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2385 = 6'h27 == _myNewVec_28_T_3[5:0] ? myVec_39 : _GEN_2384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2386 = 6'h28 == _myNewVec_28_T_3[5:0] ? myVec_40 : _GEN_2385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2387 = 6'h29 == _myNewVec_28_T_3[5:0] ? myVec_41 : _GEN_2386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2388 = 6'h2a == _myNewVec_28_T_3[5:0] ? myVec_42 : _GEN_2387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2389 = 6'h2b == _myNewVec_28_T_3[5:0] ? myVec_43 : _GEN_2388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2390 = 6'h2c == _myNewVec_28_T_3[5:0] ? myVec_44 : _GEN_2389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2391 = 6'h2d == _myNewVec_28_T_3[5:0] ? myVec_45 : _GEN_2390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2392 = 6'h2e == _myNewVec_28_T_3[5:0] ? myVec_46 : _GEN_2391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2393 = 6'h2f == _myNewVec_28_T_3[5:0] ? myVec_47 : _GEN_2392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2394 = 6'h30 == _myNewVec_28_T_3[5:0] ? myVec_48 : _GEN_2393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2395 = 6'h31 == _myNewVec_28_T_3[5:0] ? myVec_49 : _GEN_2394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2396 = 6'h32 == _myNewVec_28_T_3[5:0] ? myVec_50 : _GEN_2395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2397 = 6'h33 == _myNewVec_28_T_3[5:0] ? myVec_51 : _GEN_2396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2398 = 6'h34 == _myNewVec_28_T_3[5:0] ? myVec_52 : _GEN_2397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2399 = 6'h35 == _myNewVec_28_T_3[5:0] ? myVec_53 : _GEN_2398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2400 = 6'h36 == _myNewVec_28_T_3[5:0] ? myVec_54 : _GEN_2399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2401 = 6'h37 == _myNewVec_28_T_3[5:0] ? myVec_55 : _GEN_2400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2402 = 6'h38 == _myNewVec_28_T_3[5:0] ? myVec_56 : _GEN_2401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2403 = 6'h39 == _myNewVec_28_T_3[5:0] ? myVec_57 : _GEN_2402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2404 = 6'h3a == _myNewVec_28_T_3[5:0] ? myVec_58 : _GEN_2403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2405 = 6'h3b == _myNewVec_28_T_3[5:0] ? myVec_59 : _GEN_2404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2406 = 6'h3c == _myNewVec_28_T_3[5:0] ? myVec_60 : _GEN_2405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2407 = 6'h3d == _myNewVec_28_T_3[5:0] ? myVec_61 : _GEN_2406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2408 = 6'h3e == _myNewVec_28_T_3[5:0] ? myVec_62 : _GEN_2407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_28 = 6'h3f == _myNewVec_28_T_3[5:0] ? myVec_63 : _GEN_2408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_27_T_3 = _myNewVec_63_T_1 + 16'h24; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2411 = 6'h1 == _myNewVec_27_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2412 = 6'h2 == _myNewVec_27_T_3[5:0] ? myVec_2 : _GEN_2411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2413 = 6'h3 == _myNewVec_27_T_3[5:0] ? myVec_3 : _GEN_2412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2414 = 6'h4 == _myNewVec_27_T_3[5:0] ? myVec_4 : _GEN_2413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2415 = 6'h5 == _myNewVec_27_T_3[5:0] ? myVec_5 : _GEN_2414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2416 = 6'h6 == _myNewVec_27_T_3[5:0] ? myVec_6 : _GEN_2415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2417 = 6'h7 == _myNewVec_27_T_3[5:0] ? myVec_7 : _GEN_2416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2418 = 6'h8 == _myNewVec_27_T_3[5:0] ? myVec_8 : _GEN_2417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2419 = 6'h9 == _myNewVec_27_T_3[5:0] ? myVec_9 : _GEN_2418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2420 = 6'ha == _myNewVec_27_T_3[5:0] ? myVec_10 : _GEN_2419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2421 = 6'hb == _myNewVec_27_T_3[5:0] ? myVec_11 : _GEN_2420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2422 = 6'hc == _myNewVec_27_T_3[5:0] ? myVec_12 : _GEN_2421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2423 = 6'hd == _myNewVec_27_T_3[5:0] ? myVec_13 : _GEN_2422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2424 = 6'he == _myNewVec_27_T_3[5:0] ? myVec_14 : _GEN_2423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2425 = 6'hf == _myNewVec_27_T_3[5:0] ? myVec_15 : _GEN_2424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2426 = 6'h10 == _myNewVec_27_T_3[5:0] ? myVec_16 : _GEN_2425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2427 = 6'h11 == _myNewVec_27_T_3[5:0] ? myVec_17 : _GEN_2426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2428 = 6'h12 == _myNewVec_27_T_3[5:0] ? myVec_18 : _GEN_2427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2429 = 6'h13 == _myNewVec_27_T_3[5:0] ? myVec_19 : _GEN_2428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2430 = 6'h14 == _myNewVec_27_T_3[5:0] ? myVec_20 : _GEN_2429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2431 = 6'h15 == _myNewVec_27_T_3[5:0] ? myVec_21 : _GEN_2430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2432 = 6'h16 == _myNewVec_27_T_3[5:0] ? myVec_22 : _GEN_2431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2433 = 6'h17 == _myNewVec_27_T_3[5:0] ? myVec_23 : _GEN_2432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2434 = 6'h18 == _myNewVec_27_T_3[5:0] ? myVec_24 : _GEN_2433; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2435 = 6'h19 == _myNewVec_27_T_3[5:0] ? myVec_25 : _GEN_2434; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2436 = 6'h1a == _myNewVec_27_T_3[5:0] ? myVec_26 : _GEN_2435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2437 = 6'h1b == _myNewVec_27_T_3[5:0] ? myVec_27 : _GEN_2436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2438 = 6'h1c == _myNewVec_27_T_3[5:0] ? myVec_28 : _GEN_2437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2439 = 6'h1d == _myNewVec_27_T_3[5:0] ? myVec_29 : _GEN_2438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2440 = 6'h1e == _myNewVec_27_T_3[5:0] ? myVec_30 : _GEN_2439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2441 = 6'h1f == _myNewVec_27_T_3[5:0] ? myVec_31 : _GEN_2440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2442 = 6'h20 == _myNewVec_27_T_3[5:0] ? myVec_32 : _GEN_2441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2443 = 6'h21 == _myNewVec_27_T_3[5:0] ? myVec_33 : _GEN_2442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2444 = 6'h22 == _myNewVec_27_T_3[5:0] ? myVec_34 : _GEN_2443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2445 = 6'h23 == _myNewVec_27_T_3[5:0] ? myVec_35 : _GEN_2444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2446 = 6'h24 == _myNewVec_27_T_3[5:0] ? myVec_36 : _GEN_2445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2447 = 6'h25 == _myNewVec_27_T_3[5:0] ? myVec_37 : _GEN_2446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2448 = 6'h26 == _myNewVec_27_T_3[5:0] ? myVec_38 : _GEN_2447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2449 = 6'h27 == _myNewVec_27_T_3[5:0] ? myVec_39 : _GEN_2448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2450 = 6'h28 == _myNewVec_27_T_3[5:0] ? myVec_40 : _GEN_2449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2451 = 6'h29 == _myNewVec_27_T_3[5:0] ? myVec_41 : _GEN_2450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2452 = 6'h2a == _myNewVec_27_T_3[5:0] ? myVec_42 : _GEN_2451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2453 = 6'h2b == _myNewVec_27_T_3[5:0] ? myVec_43 : _GEN_2452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2454 = 6'h2c == _myNewVec_27_T_3[5:0] ? myVec_44 : _GEN_2453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2455 = 6'h2d == _myNewVec_27_T_3[5:0] ? myVec_45 : _GEN_2454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2456 = 6'h2e == _myNewVec_27_T_3[5:0] ? myVec_46 : _GEN_2455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2457 = 6'h2f == _myNewVec_27_T_3[5:0] ? myVec_47 : _GEN_2456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2458 = 6'h30 == _myNewVec_27_T_3[5:0] ? myVec_48 : _GEN_2457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2459 = 6'h31 == _myNewVec_27_T_3[5:0] ? myVec_49 : _GEN_2458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2460 = 6'h32 == _myNewVec_27_T_3[5:0] ? myVec_50 : _GEN_2459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2461 = 6'h33 == _myNewVec_27_T_3[5:0] ? myVec_51 : _GEN_2460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2462 = 6'h34 == _myNewVec_27_T_3[5:0] ? myVec_52 : _GEN_2461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2463 = 6'h35 == _myNewVec_27_T_3[5:0] ? myVec_53 : _GEN_2462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2464 = 6'h36 == _myNewVec_27_T_3[5:0] ? myVec_54 : _GEN_2463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2465 = 6'h37 == _myNewVec_27_T_3[5:0] ? myVec_55 : _GEN_2464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2466 = 6'h38 == _myNewVec_27_T_3[5:0] ? myVec_56 : _GEN_2465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2467 = 6'h39 == _myNewVec_27_T_3[5:0] ? myVec_57 : _GEN_2466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2468 = 6'h3a == _myNewVec_27_T_3[5:0] ? myVec_58 : _GEN_2467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2469 = 6'h3b == _myNewVec_27_T_3[5:0] ? myVec_59 : _GEN_2468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2470 = 6'h3c == _myNewVec_27_T_3[5:0] ? myVec_60 : _GEN_2469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2471 = 6'h3d == _myNewVec_27_T_3[5:0] ? myVec_61 : _GEN_2470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2472 = 6'h3e == _myNewVec_27_T_3[5:0] ? myVec_62 : _GEN_2471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_27 = 6'h3f == _myNewVec_27_T_3[5:0] ? myVec_63 : _GEN_2472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_26_T_3 = _myNewVec_63_T_1 + 16'h25; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2475 = 6'h1 == _myNewVec_26_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2476 = 6'h2 == _myNewVec_26_T_3[5:0] ? myVec_2 : _GEN_2475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2477 = 6'h3 == _myNewVec_26_T_3[5:0] ? myVec_3 : _GEN_2476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2478 = 6'h4 == _myNewVec_26_T_3[5:0] ? myVec_4 : _GEN_2477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2479 = 6'h5 == _myNewVec_26_T_3[5:0] ? myVec_5 : _GEN_2478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2480 = 6'h6 == _myNewVec_26_T_3[5:0] ? myVec_6 : _GEN_2479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2481 = 6'h7 == _myNewVec_26_T_3[5:0] ? myVec_7 : _GEN_2480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2482 = 6'h8 == _myNewVec_26_T_3[5:0] ? myVec_8 : _GEN_2481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2483 = 6'h9 == _myNewVec_26_T_3[5:0] ? myVec_9 : _GEN_2482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2484 = 6'ha == _myNewVec_26_T_3[5:0] ? myVec_10 : _GEN_2483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2485 = 6'hb == _myNewVec_26_T_3[5:0] ? myVec_11 : _GEN_2484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2486 = 6'hc == _myNewVec_26_T_3[5:0] ? myVec_12 : _GEN_2485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2487 = 6'hd == _myNewVec_26_T_3[5:0] ? myVec_13 : _GEN_2486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2488 = 6'he == _myNewVec_26_T_3[5:0] ? myVec_14 : _GEN_2487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2489 = 6'hf == _myNewVec_26_T_3[5:0] ? myVec_15 : _GEN_2488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2490 = 6'h10 == _myNewVec_26_T_3[5:0] ? myVec_16 : _GEN_2489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2491 = 6'h11 == _myNewVec_26_T_3[5:0] ? myVec_17 : _GEN_2490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2492 = 6'h12 == _myNewVec_26_T_3[5:0] ? myVec_18 : _GEN_2491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2493 = 6'h13 == _myNewVec_26_T_3[5:0] ? myVec_19 : _GEN_2492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2494 = 6'h14 == _myNewVec_26_T_3[5:0] ? myVec_20 : _GEN_2493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2495 = 6'h15 == _myNewVec_26_T_3[5:0] ? myVec_21 : _GEN_2494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2496 = 6'h16 == _myNewVec_26_T_3[5:0] ? myVec_22 : _GEN_2495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2497 = 6'h17 == _myNewVec_26_T_3[5:0] ? myVec_23 : _GEN_2496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2498 = 6'h18 == _myNewVec_26_T_3[5:0] ? myVec_24 : _GEN_2497; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2499 = 6'h19 == _myNewVec_26_T_3[5:0] ? myVec_25 : _GEN_2498; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2500 = 6'h1a == _myNewVec_26_T_3[5:0] ? myVec_26 : _GEN_2499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2501 = 6'h1b == _myNewVec_26_T_3[5:0] ? myVec_27 : _GEN_2500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2502 = 6'h1c == _myNewVec_26_T_3[5:0] ? myVec_28 : _GEN_2501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2503 = 6'h1d == _myNewVec_26_T_3[5:0] ? myVec_29 : _GEN_2502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2504 = 6'h1e == _myNewVec_26_T_3[5:0] ? myVec_30 : _GEN_2503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2505 = 6'h1f == _myNewVec_26_T_3[5:0] ? myVec_31 : _GEN_2504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2506 = 6'h20 == _myNewVec_26_T_3[5:0] ? myVec_32 : _GEN_2505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2507 = 6'h21 == _myNewVec_26_T_3[5:0] ? myVec_33 : _GEN_2506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2508 = 6'h22 == _myNewVec_26_T_3[5:0] ? myVec_34 : _GEN_2507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2509 = 6'h23 == _myNewVec_26_T_3[5:0] ? myVec_35 : _GEN_2508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2510 = 6'h24 == _myNewVec_26_T_3[5:0] ? myVec_36 : _GEN_2509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2511 = 6'h25 == _myNewVec_26_T_3[5:0] ? myVec_37 : _GEN_2510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2512 = 6'h26 == _myNewVec_26_T_3[5:0] ? myVec_38 : _GEN_2511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2513 = 6'h27 == _myNewVec_26_T_3[5:0] ? myVec_39 : _GEN_2512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2514 = 6'h28 == _myNewVec_26_T_3[5:0] ? myVec_40 : _GEN_2513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2515 = 6'h29 == _myNewVec_26_T_3[5:0] ? myVec_41 : _GEN_2514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2516 = 6'h2a == _myNewVec_26_T_3[5:0] ? myVec_42 : _GEN_2515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2517 = 6'h2b == _myNewVec_26_T_3[5:0] ? myVec_43 : _GEN_2516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2518 = 6'h2c == _myNewVec_26_T_3[5:0] ? myVec_44 : _GEN_2517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2519 = 6'h2d == _myNewVec_26_T_3[5:0] ? myVec_45 : _GEN_2518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2520 = 6'h2e == _myNewVec_26_T_3[5:0] ? myVec_46 : _GEN_2519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2521 = 6'h2f == _myNewVec_26_T_3[5:0] ? myVec_47 : _GEN_2520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2522 = 6'h30 == _myNewVec_26_T_3[5:0] ? myVec_48 : _GEN_2521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2523 = 6'h31 == _myNewVec_26_T_3[5:0] ? myVec_49 : _GEN_2522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2524 = 6'h32 == _myNewVec_26_T_3[5:0] ? myVec_50 : _GEN_2523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2525 = 6'h33 == _myNewVec_26_T_3[5:0] ? myVec_51 : _GEN_2524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2526 = 6'h34 == _myNewVec_26_T_3[5:0] ? myVec_52 : _GEN_2525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2527 = 6'h35 == _myNewVec_26_T_3[5:0] ? myVec_53 : _GEN_2526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2528 = 6'h36 == _myNewVec_26_T_3[5:0] ? myVec_54 : _GEN_2527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2529 = 6'h37 == _myNewVec_26_T_3[5:0] ? myVec_55 : _GEN_2528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2530 = 6'h38 == _myNewVec_26_T_3[5:0] ? myVec_56 : _GEN_2529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2531 = 6'h39 == _myNewVec_26_T_3[5:0] ? myVec_57 : _GEN_2530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2532 = 6'h3a == _myNewVec_26_T_3[5:0] ? myVec_58 : _GEN_2531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2533 = 6'h3b == _myNewVec_26_T_3[5:0] ? myVec_59 : _GEN_2532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2534 = 6'h3c == _myNewVec_26_T_3[5:0] ? myVec_60 : _GEN_2533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2535 = 6'h3d == _myNewVec_26_T_3[5:0] ? myVec_61 : _GEN_2534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2536 = 6'h3e == _myNewVec_26_T_3[5:0] ? myVec_62 : _GEN_2535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_26 = 6'h3f == _myNewVec_26_T_3[5:0] ? myVec_63 : _GEN_2536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_25_T_3 = _myNewVec_63_T_1 + 16'h26; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2539 = 6'h1 == _myNewVec_25_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2540 = 6'h2 == _myNewVec_25_T_3[5:0] ? myVec_2 : _GEN_2539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2541 = 6'h3 == _myNewVec_25_T_3[5:0] ? myVec_3 : _GEN_2540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2542 = 6'h4 == _myNewVec_25_T_3[5:0] ? myVec_4 : _GEN_2541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2543 = 6'h5 == _myNewVec_25_T_3[5:0] ? myVec_5 : _GEN_2542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2544 = 6'h6 == _myNewVec_25_T_3[5:0] ? myVec_6 : _GEN_2543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2545 = 6'h7 == _myNewVec_25_T_3[5:0] ? myVec_7 : _GEN_2544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2546 = 6'h8 == _myNewVec_25_T_3[5:0] ? myVec_8 : _GEN_2545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2547 = 6'h9 == _myNewVec_25_T_3[5:0] ? myVec_9 : _GEN_2546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2548 = 6'ha == _myNewVec_25_T_3[5:0] ? myVec_10 : _GEN_2547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2549 = 6'hb == _myNewVec_25_T_3[5:0] ? myVec_11 : _GEN_2548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2550 = 6'hc == _myNewVec_25_T_3[5:0] ? myVec_12 : _GEN_2549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2551 = 6'hd == _myNewVec_25_T_3[5:0] ? myVec_13 : _GEN_2550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2552 = 6'he == _myNewVec_25_T_3[5:0] ? myVec_14 : _GEN_2551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2553 = 6'hf == _myNewVec_25_T_3[5:0] ? myVec_15 : _GEN_2552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2554 = 6'h10 == _myNewVec_25_T_3[5:0] ? myVec_16 : _GEN_2553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2555 = 6'h11 == _myNewVec_25_T_3[5:0] ? myVec_17 : _GEN_2554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2556 = 6'h12 == _myNewVec_25_T_3[5:0] ? myVec_18 : _GEN_2555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2557 = 6'h13 == _myNewVec_25_T_3[5:0] ? myVec_19 : _GEN_2556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2558 = 6'h14 == _myNewVec_25_T_3[5:0] ? myVec_20 : _GEN_2557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2559 = 6'h15 == _myNewVec_25_T_3[5:0] ? myVec_21 : _GEN_2558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2560 = 6'h16 == _myNewVec_25_T_3[5:0] ? myVec_22 : _GEN_2559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2561 = 6'h17 == _myNewVec_25_T_3[5:0] ? myVec_23 : _GEN_2560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2562 = 6'h18 == _myNewVec_25_T_3[5:0] ? myVec_24 : _GEN_2561; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2563 = 6'h19 == _myNewVec_25_T_3[5:0] ? myVec_25 : _GEN_2562; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2564 = 6'h1a == _myNewVec_25_T_3[5:0] ? myVec_26 : _GEN_2563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2565 = 6'h1b == _myNewVec_25_T_3[5:0] ? myVec_27 : _GEN_2564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2566 = 6'h1c == _myNewVec_25_T_3[5:0] ? myVec_28 : _GEN_2565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2567 = 6'h1d == _myNewVec_25_T_3[5:0] ? myVec_29 : _GEN_2566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2568 = 6'h1e == _myNewVec_25_T_3[5:0] ? myVec_30 : _GEN_2567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2569 = 6'h1f == _myNewVec_25_T_3[5:0] ? myVec_31 : _GEN_2568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2570 = 6'h20 == _myNewVec_25_T_3[5:0] ? myVec_32 : _GEN_2569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2571 = 6'h21 == _myNewVec_25_T_3[5:0] ? myVec_33 : _GEN_2570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2572 = 6'h22 == _myNewVec_25_T_3[5:0] ? myVec_34 : _GEN_2571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2573 = 6'h23 == _myNewVec_25_T_3[5:0] ? myVec_35 : _GEN_2572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2574 = 6'h24 == _myNewVec_25_T_3[5:0] ? myVec_36 : _GEN_2573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2575 = 6'h25 == _myNewVec_25_T_3[5:0] ? myVec_37 : _GEN_2574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2576 = 6'h26 == _myNewVec_25_T_3[5:0] ? myVec_38 : _GEN_2575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2577 = 6'h27 == _myNewVec_25_T_3[5:0] ? myVec_39 : _GEN_2576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2578 = 6'h28 == _myNewVec_25_T_3[5:0] ? myVec_40 : _GEN_2577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2579 = 6'h29 == _myNewVec_25_T_3[5:0] ? myVec_41 : _GEN_2578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2580 = 6'h2a == _myNewVec_25_T_3[5:0] ? myVec_42 : _GEN_2579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2581 = 6'h2b == _myNewVec_25_T_3[5:0] ? myVec_43 : _GEN_2580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2582 = 6'h2c == _myNewVec_25_T_3[5:0] ? myVec_44 : _GEN_2581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2583 = 6'h2d == _myNewVec_25_T_3[5:0] ? myVec_45 : _GEN_2582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2584 = 6'h2e == _myNewVec_25_T_3[5:0] ? myVec_46 : _GEN_2583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2585 = 6'h2f == _myNewVec_25_T_3[5:0] ? myVec_47 : _GEN_2584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2586 = 6'h30 == _myNewVec_25_T_3[5:0] ? myVec_48 : _GEN_2585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2587 = 6'h31 == _myNewVec_25_T_3[5:0] ? myVec_49 : _GEN_2586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2588 = 6'h32 == _myNewVec_25_T_3[5:0] ? myVec_50 : _GEN_2587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2589 = 6'h33 == _myNewVec_25_T_3[5:0] ? myVec_51 : _GEN_2588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2590 = 6'h34 == _myNewVec_25_T_3[5:0] ? myVec_52 : _GEN_2589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2591 = 6'h35 == _myNewVec_25_T_3[5:0] ? myVec_53 : _GEN_2590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2592 = 6'h36 == _myNewVec_25_T_3[5:0] ? myVec_54 : _GEN_2591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2593 = 6'h37 == _myNewVec_25_T_3[5:0] ? myVec_55 : _GEN_2592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2594 = 6'h38 == _myNewVec_25_T_3[5:0] ? myVec_56 : _GEN_2593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2595 = 6'h39 == _myNewVec_25_T_3[5:0] ? myVec_57 : _GEN_2594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2596 = 6'h3a == _myNewVec_25_T_3[5:0] ? myVec_58 : _GEN_2595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2597 = 6'h3b == _myNewVec_25_T_3[5:0] ? myVec_59 : _GEN_2596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2598 = 6'h3c == _myNewVec_25_T_3[5:0] ? myVec_60 : _GEN_2597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2599 = 6'h3d == _myNewVec_25_T_3[5:0] ? myVec_61 : _GEN_2598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2600 = 6'h3e == _myNewVec_25_T_3[5:0] ? myVec_62 : _GEN_2599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_25 = 6'h3f == _myNewVec_25_T_3[5:0] ? myVec_63 : _GEN_2600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_24_T_3 = _myNewVec_63_T_1 + 16'h27; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2603 = 6'h1 == _myNewVec_24_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2604 = 6'h2 == _myNewVec_24_T_3[5:0] ? myVec_2 : _GEN_2603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2605 = 6'h3 == _myNewVec_24_T_3[5:0] ? myVec_3 : _GEN_2604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2606 = 6'h4 == _myNewVec_24_T_3[5:0] ? myVec_4 : _GEN_2605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2607 = 6'h5 == _myNewVec_24_T_3[5:0] ? myVec_5 : _GEN_2606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2608 = 6'h6 == _myNewVec_24_T_3[5:0] ? myVec_6 : _GEN_2607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2609 = 6'h7 == _myNewVec_24_T_3[5:0] ? myVec_7 : _GEN_2608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2610 = 6'h8 == _myNewVec_24_T_3[5:0] ? myVec_8 : _GEN_2609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2611 = 6'h9 == _myNewVec_24_T_3[5:0] ? myVec_9 : _GEN_2610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2612 = 6'ha == _myNewVec_24_T_3[5:0] ? myVec_10 : _GEN_2611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2613 = 6'hb == _myNewVec_24_T_3[5:0] ? myVec_11 : _GEN_2612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2614 = 6'hc == _myNewVec_24_T_3[5:0] ? myVec_12 : _GEN_2613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2615 = 6'hd == _myNewVec_24_T_3[5:0] ? myVec_13 : _GEN_2614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2616 = 6'he == _myNewVec_24_T_3[5:0] ? myVec_14 : _GEN_2615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2617 = 6'hf == _myNewVec_24_T_3[5:0] ? myVec_15 : _GEN_2616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2618 = 6'h10 == _myNewVec_24_T_3[5:0] ? myVec_16 : _GEN_2617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2619 = 6'h11 == _myNewVec_24_T_3[5:0] ? myVec_17 : _GEN_2618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2620 = 6'h12 == _myNewVec_24_T_3[5:0] ? myVec_18 : _GEN_2619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2621 = 6'h13 == _myNewVec_24_T_3[5:0] ? myVec_19 : _GEN_2620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2622 = 6'h14 == _myNewVec_24_T_3[5:0] ? myVec_20 : _GEN_2621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2623 = 6'h15 == _myNewVec_24_T_3[5:0] ? myVec_21 : _GEN_2622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2624 = 6'h16 == _myNewVec_24_T_3[5:0] ? myVec_22 : _GEN_2623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2625 = 6'h17 == _myNewVec_24_T_3[5:0] ? myVec_23 : _GEN_2624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2626 = 6'h18 == _myNewVec_24_T_3[5:0] ? myVec_24 : _GEN_2625; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2627 = 6'h19 == _myNewVec_24_T_3[5:0] ? myVec_25 : _GEN_2626; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2628 = 6'h1a == _myNewVec_24_T_3[5:0] ? myVec_26 : _GEN_2627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2629 = 6'h1b == _myNewVec_24_T_3[5:0] ? myVec_27 : _GEN_2628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2630 = 6'h1c == _myNewVec_24_T_3[5:0] ? myVec_28 : _GEN_2629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2631 = 6'h1d == _myNewVec_24_T_3[5:0] ? myVec_29 : _GEN_2630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2632 = 6'h1e == _myNewVec_24_T_3[5:0] ? myVec_30 : _GEN_2631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2633 = 6'h1f == _myNewVec_24_T_3[5:0] ? myVec_31 : _GEN_2632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2634 = 6'h20 == _myNewVec_24_T_3[5:0] ? myVec_32 : _GEN_2633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2635 = 6'h21 == _myNewVec_24_T_3[5:0] ? myVec_33 : _GEN_2634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2636 = 6'h22 == _myNewVec_24_T_3[5:0] ? myVec_34 : _GEN_2635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2637 = 6'h23 == _myNewVec_24_T_3[5:0] ? myVec_35 : _GEN_2636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2638 = 6'h24 == _myNewVec_24_T_3[5:0] ? myVec_36 : _GEN_2637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2639 = 6'h25 == _myNewVec_24_T_3[5:0] ? myVec_37 : _GEN_2638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2640 = 6'h26 == _myNewVec_24_T_3[5:0] ? myVec_38 : _GEN_2639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2641 = 6'h27 == _myNewVec_24_T_3[5:0] ? myVec_39 : _GEN_2640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2642 = 6'h28 == _myNewVec_24_T_3[5:0] ? myVec_40 : _GEN_2641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2643 = 6'h29 == _myNewVec_24_T_3[5:0] ? myVec_41 : _GEN_2642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2644 = 6'h2a == _myNewVec_24_T_3[5:0] ? myVec_42 : _GEN_2643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2645 = 6'h2b == _myNewVec_24_T_3[5:0] ? myVec_43 : _GEN_2644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2646 = 6'h2c == _myNewVec_24_T_3[5:0] ? myVec_44 : _GEN_2645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2647 = 6'h2d == _myNewVec_24_T_3[5:0] ? myVec_45 : _GEN_2646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2648 = 6'h2e == _myNewVec_24_T_3[5:0] ? myVec_46 : _GEN_2647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2649 = 6'h2f == _myNewVec_24_T_3[5:0] ? myVec_47 : _GEN_2648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2650 = 6'h30 == _myNewVec_24_T_3[5:0] ? myVec_48 : _GEN_2649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2651 = 6'h31 == _myNewVec_24_T_3[5:0] ? myVec_49 : _GEN_2650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2652 = 6'h32 == _myNewVec_24_T_3[5:0] ? myVec_50 : _GEN_2651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2653 = 6'h33 == _myNewVec_24_T_3[5:0] ? myVec_51 : _GEN_2652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2654 = 6'h34 == _myNewVec_24_T_3[5:0] ? myVec_52 : _GEN_2653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2655 = 6'h35 == _myNewVec_24_T_3[5:0] ? myVec_53 : _GEN_2654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2656 = 6'h36 == _myNewVec_24_T_3[5:0] ? myVec_54 : _GEN_2655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2657 = 6'h37 == _myNewVec_24_T_3[5:0] ? myVec_55 : _GEN_2656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2658 = 6'h38 == _myNewVec_24_T_3[5:0] ? myVec_56 : _GEN_2657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2659 = 6'h39 == _myNewVec_24_T_3[5:0] ? myVec_57 : _GEN_2658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2660 = 6'h3a == _myNewVec_24_T_3[5:0] ? myVec_58 : _GEN_2659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2661 = 6'h3b == _myNewVec_24_T_3[5:0] ? myVec_59 : _GEN_2660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2662 = 6'h3c == _myNewVec_24_T_3[5:0] ? myVec_60 : _GEN_2661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2663 = 6'h3d == _myNewVec_24_T_3[5:0] ? myVec_61 : _GEN_2662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2664 = 6'h3e == _myNewVec_24_T_3[5:0] ? myVec_62 : _GEN_2663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_24 = 6'h3f == _myNewVec_24_T_3[5:0] ? myVec_63 : _GEN_2664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_23_T_3 = _myNewVec_63_T_1 + 16'h28; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2667 = 6'h1 == _myNewVec_23_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2668 = 6'h2 == _myNewVec_23_T_3[5:0] ? myVec_2 : _GEN_2667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2669 = 6'h3 == _myNewVec_23_T_3[5:0] ? myVec_3 : _GEN_2668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2670 = 6'h4 == _myNewVec_23_T_3[5:0] ? myVec_4 : _GEN_2669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2671 = 6'h5 == _myNewVec_23_T_3[5:0] ? myVec_5 : _GEN_2670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2672 = 6'h6 == _myNewVec_23_T_3[5:0] ? myVec_6 : _GEN_2671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2673 = 6'h7 == _myNewVec_23_T_3[5:0] ? myVec_7 : _GEN_2672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2674 = 6'h8 == _myNewVec_23_T_3[5:0] ? myVec_8 : _GEN_2673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2675 = 6'h9 == _myNewVec_23_T_3[5:0] ? myVec_9 : _GEN_2674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2676 = 6'ha == _myNewVec_23_T_3[5:0] ? myVec_10 : _GEN_2675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2677 = 6'hb == _myNewVec_23_T_3[5:0] ? myVec_11 : _GEN_2676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2678 = 6'hc == _myNewVec_23_T_3[5:0] ? myVec_12 : _GEN_2677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2679 = 6'hd == _myNewVec_23_T_3[5:0] ? myVec_13 : _GEN_2678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2680 = 6'he == _myNewVec_23_T_3[5:0] ? myVec_14 : _GEN_2679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2681 = 6'hf == _myNewVec_23_T_3[5:0] ? myVec_15 : _GEN_2680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2682 = 6'h10 == _myNewVec_23_T_3[5:0] ? myVec_16 : _GEN_2681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2683 = 6'h11 == _myNewVec_23_T_3[5:0] ? myVec_17 : _GEN_2682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2684 = 6'h12 == _myNewVec_23_T_3[5:0] ? myVec_18 : _GEN_2683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2685 = 6'h13 == _myNewVec_23_T_3[5:0] ? myVec_19 : _GEN_2684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2686 = 6'h14 == _myNewVec_23_T_3[5:0] ? myVec_20 : _GEN_2685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2687 = 6'h15 == _myNewVec_23_T_3[5:0] ? myVec_21 : _GEN_2686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2688 = 6'h16 == _myNewVec_23_T_3[5:0] ? myVec_22 : _GEN_2687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2689 = 6'h17 == _myNewVec_23_T_3[5:0] ? myVec_23 : _GEN_2688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2690 = 6'h18 == _myNewVec_23_T_3[5:0] ? myVec_24 : _GEN_2689; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2691 = 6'h19 == _myNewVec_23_T_3[5:0] ? myVec_25 : _GEN_2690; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2692 = 6'h1a == _myNewVec_23_T_3[5:0] ? myVec_26 : _GEN_2691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2693 = 6'h1b == _myNewVec_23_T_3[5:0] ? myVec_27 : _GEN_2692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2694 = 6'h1c == _myNewVec_23_T_3[5:0] ? myVec_28 : _GEN_2693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2695 = 6'h1d == _myNewVec_23_T_3[5:0] ? myVec_29 : _GEN_2694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2696 = 6'h1e == _myNewVec_23_T_3[5:0] ? myVec_30 : _GEN_2695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2697 = 6'h1f == _myNewVec_23_T_3[5:0] ? myVec_31 : _GEN_2696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2698 = 6'h20 == _myNewVec_23_T_3[5:0] ? myVec_32 : _GEN_2697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2699 = 6'h21 == _myNewVec_23_T_3[5:0] ? myVec_33 : _GEN_2698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2700 = 6'h22 == _myNewVec_23_T_3[5:0] ? myVec_34 : _GEN_2699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2701 = 6'h23 == _myNewVec_23_T_3[5:0] ? myVec_35 : _GEN_2700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2702 = 6'h24 == _myNewVec_23_T_3[5:0] ? myVec_36 : _GEN_2701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2703 = 6'h25 == _myNewVec_23_T_3[5:0] ? myVec_37 : _GEN_2702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2704 = 6'h26 == _myNewVec_23_T_3[5:0] ? myVec_38 : _GEN_2703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2705 = 6'h27 == _myNewVec_23_T_3[5:0] ? myVec_39 : _GEN_2704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2706 = 6'h28 == _myNewVec_23_T_3[5:0] ? myVec_40 : _GEN_2705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2707 = 6'h29 == _myNewVec_23_T_3[5:0] ? myVec_41 : _GEN_2706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2708 = 6'h2a == _myNewVec_23_T_3[5:0] ? myVec_42 : _GEN_2707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2709 = 6'h2b == _myNewVec_23_T_3[5:0] ? myVec_43 : _GEN_2708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2710 = 6'h2c == _myNewVec_23_T_3[5:0] ? myVec_44 : _GEN_2709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2711 = 6'h2d == _myNewVec_23_T_3[5:0] ? myVec_45 : _GEN_2710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2712 = 6'h2e == _myNewVec_23_T_3[5:0] ? myVec_46 : _GEN_2711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2713 = 6'h2f == _myNewVec_23_T_3[5:0] ? myVec_47 : _GEN_2712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2714 = 6'h30 == _myNewVec_23_T_3[5:0] ? myVec_48 : _GEN_2713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2715 = 6'h31 == _myNewVec_23_T_3[5:0] ? myVec_49 : _GEN_2714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2716 = 6'h32 == _myNewVec_23_T_3[5:0] ? myVec_50 : _GEN_2715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2717 = 6'h33 == _myNewVec_23_T_3[5:0] ? myVec_51 : _GEN_2716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2718 = 6'h34 == _myNewVec_23_T_3[5:0] ? myVec_52 : _GEN_2717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2719 = 6'h35 == _myNewVec_23_T_3[5:0] ? myVec_53 : _GEN_2718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2720 = 6'h36 == _myNewVec_23_T_3[5:0] ? myVec_54 : _GEN_2719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2721 = 6'h37 == _myNewVec_23_T_3[5:0] ? myVec_55 : _GEN_2720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2722 = 6'h38 == _myNewVec_23_T_3[5:0] ? myVec_56 : _GEN_2721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2723 = 6'h39 == _myNewVec_23_T_3[5:0] ? myVec_57 : _GEN_2722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2724 = 6'h3a == _myNewVec_23_T_3[5:0] ? myVec_58 : _GEN_2723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2725 = 6'h3b == _myNewVec_23_T_3[5:0] ? myVec_59 : _GEN_2724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2726 = 6'h3c == _myNewVec_23_T_3[5:0] ? myVec_60 : _GEN_2725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2727 = 6'h3d == _myNewVec_23_T_3[5:0] ? myVec_61 : _GEN_2726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2728 = 6'h3e == _myNewVec_23_T_3[5:0] ? myVec_62 : _GEN_2727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_23 = 6'h3f == _myNewVec_23_T_3[5:0] ? myVec_63 : _GEN_2728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_22_T_3 = _myNewVec_63_T_1 + 16'h29; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2731 = 6'h1 == _myNewVec_22_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2732 = 6'h2 == _myNewVec_22_T_3[5:0] ? myVec_2 : _GEN_2731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2733 = 6'h3 == _myNewVec_22_T_3[5:0] ? myVec_3 : _GEN_2732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2734 = 6'h4 == _myNewVec_22_T_3[5:0] ? myVec_4 : _GEN_2733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2735 = 6'h5 == _myNewVec_22_T_3[5:0] ? myVec_5 : _GEN_2734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2736 = 6'h6 == _myNewVec_22_T_3[5:0] ? myVec_6 : _GEN_2735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2737 = 6'h7 == _myNewVec_22_T_3[5:0] ? myVec_7 : _GEN_2736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2738 = 6'h8 == _myNewVec_22_T_3[5:0] ? myVec_8 : _GEN_2737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2739 = 6'h9 == _myNewVec_22_T_3[5:0] ? myVec_9 : _GEN_2738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2740 = 6'ha == _myNewVec_22_T_3[5:0] ? myVec_10 : _GEN_2739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2741 = 6'hb == _myNewVec_22_T_3[5:0] ? myVec_11 : _GEN_2740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2742 = 6'hc == _myNewVec_22_T_3[5:0] ? myVec_12 : _GEN_2741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2743 = 6'hd == _myNewVec_22_T_3[5:0] ? myVec_13 : _GEN_2742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2744 = 6'he == _myNewVec_22_T_3[5:0] ? myVec_14 : _GEN_2743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2745 = 6'hf == _myNewVec_22_T_3[5:0] ? myVec_15 : _GEN_2744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2746 = 6'h10 == _myNewVec_22_T_3[5:0] ? myVec_16 : _GEN_2745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2747 = 6'h11 == _myNewVec_22_T_3[5:0] ? myVec_17 : _GEN_2746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2748 = 6'h12 == _myNewVec_22_T_3[5:0] ? myVec_18 : _GEN_2747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2749 = 6'h13 == _myNewVec_22_T_3[5:0] ? myVec_19 : _GEN_2748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2750 = 6'h14 == _myNewVec_22_T_3[5:0] ? myVec_20 : _GEN_2749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2751 = 6'h15 == _myNewVec_22_T_3[5:0] ? myVec_21 : _GEN_2750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2752 = 6'h16 == _myNewVec_22_T_3[5:0] ? myVec_22 : _GEN_2751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2753 = 6'h17 == _myNewVec_22_T_3[5:0] ? myVec_23 : _GEN_2752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2754 = 6'h18 == _myNewVec_22_T_3[5:0] ? myVec_24 : _GEN_2753; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2755 = 6'h19 == _myNewVec_22_T_3[5:0] ? myVec_25 : _GEN_2754; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2756 = 6'h1a == _myNewVec_22_T_3[5:0] ? myVec_26 : _GEN_2755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2757 = 6'h1b == _myNewVec_22_T_3[5:0] ? myVec_27 : _GEN_2756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2758 = 6'h1c == _myNewVec_22_T_3[5:0] ? myVec_28 : _GEN_2757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2759 = 6'h1d == _myNewVec_22_T_3[5:0] ? myVec_29 : _GEN_2758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2760 = 6'h1e == _myNewVec_22_T_3[5:0] ? myVec_30 : _GEN_2759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2761 = 6'h1f == _myNewVec_22_T_3[5:0] ? myVec_31 : _GEN_2760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2762 = 6'h20 == _myNewVec_22_T_3[5:0] ? myVec_32 : _GEN_2761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2763 = 6'h21 == _myNewVec_22_T_3[5:0] ? myVec_33 : _GEN_2762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2764 = 6'h22 == _myNewVec_22_T_3[5:0] ? myVec_34 : _GEN_2763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2765 = 6'h23 == _myNewVec_22_T_3[5:0] ? myVec_35 : _GEN_2764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2766 = 6'h24 == _myNewVec_22_T_3[5:0] ? myVec_36 : _GEN_2765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2767 = 6'h25 == _myNewVec_22_T_3[5:0] ? myVec_37 : _GEN_2766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2768 = 6'h26 == _myNewVec_22_T_3[5:0] ? myVec_38 : _GEN_2767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2769 = 6'h27 == _myNewVec_22_T_3[5:0] ? myVec_39 : _GEN_2768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2770 = 6'h28 == _myNewVec_22_T_3[5:0] ? myVec_40 : _GEN_2769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2771 = 6'h29 == _myNewVec_22_T_3[5:0] ? myVec_41 : _GEN_2770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2772 = 6'h2a == _myNewVec_22_T_3[5:0] ? myVec_42 : _GEN_2771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2773 = 6'h2b == _myNewVec_22_T_3[5:0] ? myVec_43 : _GEN_2772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2774 = 6'h2c == _myNewVec_22_T_3[5:0] ? myVec_44 : _GEN_2773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2775 = 6'h2d == _myNewVec_22_T_3[5:0] ? myVec_45 : _GEN_2774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2776 = 6'h2e == _myNewVec_22_T_3[5:0] ? myVec_46 : _GEN_2775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2777 = 6'h2f == _myNewVec_22_T_3[5:0] ? myVec_47 : _GEN_2776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2778 = 6'h30 == _myNewVec_22_T_3[5:0] ? myVec_48 : _GEN_2777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2779 = 6'h31 == _myNewVec_22_T_3[5:0] ? myVec_49 : _GEN_2778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2780 = 6'h32 == _myNewVec_22_T_3[5:0] ? myVec_50 : _GEN_2779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2781 = 6'h33 == _myNewVec_22_T_3[5:0] ? myVec_51 : _GEN_2780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2782 = 6'h34 == _myNewVec_22_T_3[5:0] ? myVec_52 : _GEN_2781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2783 = 6'h35 == _myNewVec_22_T_3[5:0] ? myVec_53 : _GEN_2782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2784 = 6'h36 == _myNewVec_22_T_3[5:0] ? myVec_54 : _GEN_2783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2785 = 6'h37 == _myNewVec_22_T_3[5:0] ? myVec_55 : _GEN_2784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2786 = 6'h38 == _myNewVec_22_T_3[5:0] ? myVec_56 : _GEN_2785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2787 = 6'h39 == _myNewVec_22_T_3[5:0] ? myVec_57 : _GEN_2786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2788 = 6'h3a == _myNewVec_22_T_3[5:0] ? myVec_58 : _GEN_2787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2789 = 6'h3b == _myNewVec_22_T_3[5:0] ? myVec_59 : _GEN_2788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2790 = 6'h3c == _myNewVec_22_T_3[5:0] ? myVec_60 : _GEN_2789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2791 = 6'h3d == _myNewVec_22_T_3[5:0] ? myVec_61 : _GEN_2790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2792 = 6'h3e == _myNewVec_22_T_3[5:0] ? myVec_62 : _GEN_2791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_22 = 6'h3f == _myNewVec_22_T_3[5:0] ? myVec_63 : _GEN_2792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_21_T_3 = _myNewVec_63_T_1 + 16'h2a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2795 = 6'h1 == _myNewVec_21_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2796 = 6'h2 == _myNewVec_21_T_3[5:0] ? myVec_2 : _GEN_2795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2797 = 6'h3 == _myNewVec_21_T_3[5:0] ? myVec_3 : _GEN_2796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2798 = 6'h4 == _myNewVec_21_T_3[5:0] ? myVec_4 : _GEN_2797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2799 = 6'h5 == _myNewVec_21_T_3[5:0] ? myVec_5 : _GEN_2798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2800 = 6'h6 == _myNewVec_21_T_3[5:0] ? myVec_6 : _GEN_2799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2801 = 6'h7 == _myNewVec_21_T_3[5:0] ? myVec_7 : _GEN_2800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2802 = 6'h8 == _myNewVec_21_T_3[5:0] ? myVec_8 : _GEN_2801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2803 = 6'h9 == _myNewVec_21_T_3[5:0] ? myVec_9 : _GEN_2802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2804 = 6'ha == _myNewVec_21_T_3[5:0] ? myVec_10 : _GEN_2803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2805 = 6'hb == _myNewVec_21_T_3[5:0] ? myVec_11 : _GEN_2804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2806 = 6'hc == _myNewVec_21_T_3[5:0] ? myVec_12 : _GEN_2805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2807 = 6'hd == _myNewVec_21_T_3[5:0] ? myVec_13 : _GEN_2806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2808 = 6'he == _myNewVec_21_T_3[5:0] ? myVec_14 : _GEN_2807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2809 = 6'hf == _myNewVec_21_T_3[5:0] ? myVec_15 : _GEN_2808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2810 = 6'h10 == _myNewVec_21_T_3[5:0] ? myVec_16 : _GEN_2809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2811 = 6'h11 == _myNewVec_21_T_3[5:0] ? myVec_17 : _GEN_2810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2812 = 6'h12 == _myNewVec_21_T_3[5:0] ? myVec_18 : _GEN_2811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2813 = 6'h13 == _myNewVec_21_T_3[5:0] ? myVec_19 : _GEN_2812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2814 = 6'h14 == _myNewVec_21_T_3[5:0] ? myVec_20 : _GEN_2813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2815 = 6'h15 == _myNewVec_21_T_3[5:0] ? myVec_21 : _GEN_2814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2816 = 6'h16 == _myNewVec_21_T_3[5:0] ? myVec_22 : _GEN_2815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2817 = 6'h17 == _myNewVec_21_T_3[5:0] ? myVec_23 : _GEN_2816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2818 = 6'h18 == _myNewVec_21_T_3[5:0] ? myVec_24 : _GEN_2817; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2819 = 6'h19 == _myNewVec_21_T_3[5:0] ? myVec_25 : _GEN_2818; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2820 = 6'h1a == _myNewVec_21_T_3[5:0] ? myVec_26 : _GEN_2819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2821 = 6'h1b == _myNewVec_21_T_3[5:0] ? myVec_27 : _GEN_2820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2822 = 6'h1c == _myNewVec_21_T_3[5:0] ? myVec_28 : _GEN_2821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2823 = 6'h1d == _myNewVec_21_T_3[5:0] ? myVec_29 : _GEN_2822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2824 = 6'h1e == _myNewVec_21_T_3[5:0] ? myVec_30 : _GEN_2823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2825 = 6'h1f == _myNewVec_21_T_3[5:0] ? myVec_31 : _GEN_2824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2826 = 6'h20 == _myNewVec_21_T_3[5:0] ? myVec_32 : _GEN_2825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2827 = 6'h21 == _myNewVec_21_T_3[5:0] ? myVec_33 : _GEN_2826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2828 = 6'h22 == _myNewVec_21_T_3[5:0] ? myVec_34 : _GEN_2827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2829 = 6'h23 == _myNewVec_21_T_3[5:0] ? myVec_35 : _GEN_2828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2830 = 6'h24 == _myNewVec_21_T_3[5:0] ? myVec_36 : _GEN_2829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2831 = 6'h25 == _myNewVec_21_T_3[5:0] ? myVec_37 : _GEN_2830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2832 = 6'h26 == _myNewVec_21_T_3[5:0] ? myVec_38 : _GEN_2831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2833 = 6'h27 == _myNewVec_21_T_3[5:0] ? myVec_39 : _GEN_2832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2834 = 6'h28 == _myNewVec_21_T_3[5:0] ? myVec_40 : _GEN_2833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2835 = 6'h29 == _myNewVec_21_T_3[5:0] ? myVec_41 : _GEN_2834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2836 = 6'h2a == _myNewVec_21_T_3[5:0] ? myVec_42 : _GEN_2835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2837 = 6'h2b == _myNewVec_21_T_3[5:0] ? myVec_43 : _GEN_2836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2838 = 6'h2c == _myNewVec_21_T_3[5:0] ? myVec_44 : _GEN_2837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2839 = 6'h2d == _myNewVec_21_T_3[5:0] ? myVec_45 : _GEN_2838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2840 = 6'h2e == _myNewVec_21_T_3[5:0] ? myVec_46 : _GEN_2839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2841 = 6'h2f == _myNewVec_21_T_3[5:0] ? myVec_47 : _GEN_2840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2842 = 6'h30 == _myNewVec_21_T_3[5:0] ? myVec_48 : _GEN_2841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2843 = 6'h31 == _myNewVec_21_T_3[5:0] ? myVec_49 : _GEN_2842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2844 = 6'h32 == _myNewVec_21_T_3[5:0] ? myVec_50 : _GEN_2843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2845 = 6'h33 == _myNewVec_21_T_3[5:0] ? myVec_51 : _GEN_2844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2846 = 6'h34 == _myNewVec_21_T_3[5:0] ? myVec_52 : _GEN_2845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2847 = 6'h35 == _myNewVec_21_T_3[5:0] ? myVec_53 : _GEN_2846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2848 = 6'h36 == _myNewVec_21_T_3[5:0] ? myVec_54 : _GEN_2847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2849 = 6'h37 == _myNewVec_21_T_3[5:0] ? myVec_55 : _GEN_2848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2850 = 6'h38 == _myNewVec_21_T_3[5:0] ? myVec_56 : _GEN_2849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2851 = 6'h39 == _myNewVec_21_T_3[5:0] ? myVec_57 : _GEN_2850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2852 = 6'h3a == _myNewVec_21_T_3[5:0] ? myVec_58 : _GEN_2851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2853 = 6'h3b == _myNewVec_21_T_3[5:0] ? myVec_59 : _GEN_2852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2854 = 6'h3c == _myNewVec_21_T_3[5:0] ? myVec_60 : _GEN_2853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2855 = 6'h3d == _myNewVec_21_T_3[5:0] ? myVec_61 : _GEN_2854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2856 = 6'h3e == _myNewVec_21_T_3[5:0] ? myVec_62 : _GEN_2855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_21 = 6'h3f == _myNewVec_21_T_3[5:0] ? myVec_63 : _GEN_2856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_20_T_3 = _myNewVec_63_T_1 + 16'h2b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2859 = 6'h1 == _myNewVec_20_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2860 = 6'h2 == _myNewVec_20_T_3[5:0] ? myVec_2 : _GEN_2859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2861 = 6'h3 == _myNewVec_20_T_3[5:0] ? myVec_3 : _GEN_2860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2862 = 6'h4 == _myNewVec_20_T_3[5:0] ? myVec_4 : _GEN_2861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2863 = 6'h5 == _myNewVec_20_T_3[5:0] ? myVec_5 : _GEN_2862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2864 = 6'h6 == _myNewVec_20_T_3[5:0] ? myVec_6 : _GEN_2863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2865 = 6'h7 == _myNewVec_20_T_3[5:0] ? myVec_7 : _GEN_2864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2866 = 6'h8 == _myNewVec_20_T_3[5:0] ? myVec_8 : _GEN_2865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2867 = 6'h9 == _myNewVec_20_T_3[5:0] ? myVec_9 : _GEN_2866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2868 = 6'ha == _myNewVec_20_T_3[5:0] ? myVec_10 : _GEN_2867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2869 = 6'hb == _myNewVec_20_T_3[5:0] ? myVec_11 : _GEN_2868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2870 = 6'hc == _myNewVec_20_T_3[5:0] ? myVec_12 : _GEN_2869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2871 = 6'hd == _myNewVec_20_T_3[5:0] ? myVec_13 : _GEN_2870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2872 = 6'he == _myNewVec_20_T_3[5:0] ? myVec_14 : _GEN_2871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2873 = 6'hf == _myNewVec_20_T_3[5:0] ? myVec_15 : _GEN_2872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2874 = 6'h10 == _myNewVec_20_T_3[5:0] ? myVec_16 : _GEN_2873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2875 = 6'h11 == _myNewVec_20_T_3[5:0] ? myVec_17 : _GEN_2874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2876 = 6'h12 == _myNewVec_20_T_3[5:0] ? myVec_18 : _GEN_2875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2877 = 6'h13 == _myNewVec_20_T_3[5:0] ? myVec_19 : _GEN_2876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2878 = 6'h14 == _myNewVec_20_T_3[5:0] ? myVec_20 : _GEN_2877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2879 = 6'h15 == _myNewVec_20_T_3[5:0] ? myVec_21 : _GEN_2878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2880 = 6'h16 == _myNewVec_20_T_3[5:0] ? myVec_22 : _GEN_2879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2881 = 6'h17 == _myNewVec_20_T_3[5:0] ? myVec_23 : _GEN_2880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2882 = 6'h18 == _myNewVec_20_T_3[5:0] ? myVec_24 : _GEN_2881; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2883 = 6'h19 == _myNewVec_20_T_3[5:0] ? myVec_25 : _GEN_2882; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2884 = 6'h1a == _myNewVec_20_T_3[5:0] ? myVec_26 : _GEN_2883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2885 = 6'h1b == _myNewVec_20_T_3[5:0] ? myVec_27 : _GEN_2884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2886 = 6'h1c == _myNewVec_20_T_3[5:0] ? myVec_28 : _GEN_2885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2887 = 6'h1d == _myNewVec_20_T_3[5:0] ? myVec_29 : _GEN_2886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2888 = 6'h1e == _myNewVec_20_T_3[5:0] ? myVec_30 : _GEN_2887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2889 = 6'h1f == _myNewVec_20_T_3[5:0] ? myVec_31 : _GEN_2888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2890 = 6'h20 == _myNewVec_20_T_3[5:0] ? myVec_32 : _GEN_2889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2891 = 6'h21 == _myNewVec_20_T_3[5:0] ? myVec_33 : _GEN_2890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2892 = 6'h22 == _myNewVec_20_T_3[5:0] ? myVec_34 : _GEN_2891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2893 = 6'h23 == _myNewVec_20_T_3[5:0] ? myVec_35 : _GEN_2892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2894 = 6'h24 == _myNewVec_20_T_3[5:0] ? myVec_36 : _GEN_2893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2895 = 6'h25 == _myNewVec_20_T_3[5:0] ? myVec_37 : _GEN_2894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2896 = 6'h26 == _myNewVec_20_T_3[5:0] ? myVec_38 : _GEN_2895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2897 = 6'h27 == _myNewVec_20_T_3[5:0] ? myVec_39 : _GEN_2896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2898 = 6'h28 == _myNewVec_20_T_3[5:0] ? myVec_40 : _GEN_2897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2899 = 6'h29 == _myNewVec_20_T_3[5:0] ? myVec_41 : _GEN_2898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2900 = 6'h2a == _myNewVec_20_T_3[5:0] ? myVec_42 : _GEN_2899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2901 = 6'h2b == _myNewVec_20_T_3[5:0] ? myVec_43 : _GEN_2900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2902 = 6'h2c == _myNewVec_20_T_3[5:0] ? myVec_44 : _GEN_2901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2903 = 6'h2d == _myNewVec_20_T_3[5:0] ? myVec_45 : _GEN_2902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2904 = 6'h2e == _myNewVec_20_T_3[5:0] ? myVec_46 : _GEN_2903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2905 = 6'h2f == _myNewVec_20_T_3[5:0] ? myVec_47 : _GEN_2904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2906 = 6'h30 == _myNewVec_20_T_3[5:0] ? myVec_48 : _GEN_2905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2907 = 6'h31 == _myNewVec_20_T_3[5:0] ? myVec_49 : _GEN_2906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2908 = 6'h32 == _myNewVec_20_T_3[5:0] ? myVec_50 : _GEN_2907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2909 = 6'h33 == _myNewVec_20_T_3[5:0] ? myVec_51 : _GEN_2908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2910 = 6'h34 == _myNewVec_20_T_3[5:0] ? myVec_52 : _GEN_2909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2911 = 6'h35 == _myNewVec_20_T_3[5:0] ? myVec_53 : _GEN_2910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2912 = 6'h36 == _myNewVec_20_T_3[5:0] ? myVec_54 : _GEN_2911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2913 = 6'h37 == _myNewVec_20_T_3[5:0] ? myVec_55 : _GEN_2912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2914 = 6'h38 == _myNewVec_20_T_3[5:0] ? myVec_56 : _GEN_2913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2915 = 6'h39 == _myNewVec_20_T_3[5:0] ? myVec_57 : _GEN_2914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2916 = 6'h3a == _myNewVec_20_T_3[5:0] ? myVec_58 : _GEN_2915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2917 = 6'h3b == _myNewVec_20_T_3[5:0] ? myVec_59 : _GEN_2916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2918 = 6'h3c == _myNewVec_20_T_3[5:0] ? myVec_60 : _GEN_2917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2919 = 6'h3d == _myNewVec_20_T_3[5:0] ? myVec_61 : _GEN_2918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2920 = 6'h3e == _myNewVec_20_T_3[5:0] ? myVec_62 : _GEN_2919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_20 = 6'h3f == _myNewVec_20_T_3[5:0] ? myVec_63 : _GEN_2920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_19_T_3 = _myNewVec_63_T_1 + 16'h2c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2923 = 6'h1 == _myNewVec_19_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2924 = 6'h2 == _myNewVec_19_T_3[5:0] ? myVec_2 : _GEN_2923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2925 = 6'h3 == _myNewVec_19_T_3[5:0] ? myVec_3 : _GEN_2924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2926 = 6'h4 == _myNewVec_19_T_3[5:0] ? myVec_4 : _GEN_2925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2927 = 6'h5 == _myNewVec_19_T_3[5:0] ? myVec_5 : _GEN_2926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2928 = 6'h6 == _myNewVec_19_T_3[5:0] ? myVec_6 : _GEN_2927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2929 = 6'h7 == _myNewVec_19_T_3[5:0] ? myVec_7 : _GEN_2928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2930 = 6'h8 == _myNewVec_19_T_3[5:0] ? myVec_8 : _GEN_2929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2931 = 6'h9 == _myNewVec_19_T_3[5:0] ? myVec_9 : _GEN_2930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2932 = 6'ha == _myNewVec_19_T_3[5:0] ? myVec_10 : _GEN_2931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2933 = 6'hb == _myNewVec_19_T_3[5:0] ? myVec_11 : _GEN_2932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2934 = 6'hc == _myNewVec_19_T_3[5:0] ? myVec_12 : _GEN_2933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2935 = 6'hd == _myNewVec_19_T_3[5:0] ? myVec_13 : _GEN_2934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2936 = 6'he == _myNewVec_19_T_3[5:0] ? myVec_14 : _GEN_2935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2937 = 6'hf == _myNewVec_19_T_3[5:0] ? myVec_15 : _GEN_2936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2938 = 6'h10 == _myNewVec_19_T_3[5:0] ? myVec_16 : _GEN_2937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2939 = 6'h11 == _myNewVec_19_T_3[5:0] ? myVec_17 : _GEN_2938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2940 = 6'h12 == _myNewVec_19_T_3[5:0] ? myVec_18 : _GEN_2939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2941 = 6'h13 == _myNewVec_19_T_3[5:0] ? myVec_19 : _GEN_2940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2942 = 6'h14 == _myNewVec_19_T_3[5:0] ? myVec_20 : _GEN_2941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2943 = 6'h15 == _myNewVec_19_T_3[5:0] ? myVec_21 : _GEN_2942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2944 = 6'h16 == _myNewVec_19_T_3[5:0] ? myVec_22 : _GEN_2943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2945 = 6'h17 == _myNewVec_19_T_3[5:0] ? myVec_23 : _GEN_2944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2946 = 6'h18 == _myNewVec_19_T_3[5:0] ? myVec_24 : _GEN_2945; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2947 = 6'h19 == _myNewVec_19_T_3[5:0] ? myVec_25 : _GEN_2946; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2948 = 6'h1a == _myNewVec_19_T_3[5:0] ? myVec_26 : _GEN_2947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2949 = 6'h1b == _myNewVec_19_T_3[5:0] ? myVec_27 : _GEN_2948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2950 = 6'h1c == _myNewVec_19_T_3[5:0] ? myVec_28 : _GEN_2949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2951 = 6'h1d == _myNewVec_19_T_3[5:0] ? myVec_29 : _GEN_2950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2952 = 6'h1e == _myNewVec_19_T_3[5:0] ? myVec_30 : _GEN_2951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2953 = 6'h1f == _myNewVec_19_T_3[5:0] ? myVec_31 : _GEN_2952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2954 = 6'h20 == _myNewVec_19_T_3[5:0] ? myVec_32 : _GEN_2953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2955 = 6'h21 == _myNewVec_19_T_3[5:0] ? myVec_33 : _GEN_2954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2956 = 6'h22 == _myNewVec_19_T_3[5:0] ? myVec_34 : _GEN_2955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2957 = 6'h23 == _myNewVec_19_T_3[5:0] ? myVec_35 : _GEN_2956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2958 = 6'h24 == _myNewVec_19_T_3[5:0] ? myVec_36 : _GEN_2957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2959 = 6'h25 == _myNewVec_19_T_3[5:0] ? myVec_37 : _GEN_2958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2960 = 6'h26 == _myNewVec_19_T_3[5:0] ? myVec_38 : _GEN_2959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2961 = 6'h27 == _myNewVec_19_T_3[5:0] ? myVec_39 : _GEN_2960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2962 = 6'h28 == _myNewVec_19_T_3[5:0] ? myVec_40 : _GEN_2961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2963 = 6'h29 == _myNewVec_19_T_3[5:0] ? myVec_41 : _GEN_2962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2964 = 6'h2a == _myNewVec_19_T_3[5:0] ? myVec_42 : _GEN_2963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2965 = 6'h2b == _myNewVec_19_T_3[5:0] ? myVec_43 : _GEN_2964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2966 = 6'h2c == _myNewVec_19_T_3[5:0] ? myVec_44 : _GEN_2965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2967 = 6'h2d == _myNewVec_19_T_3[5:0] ? myVec_45 : _GEN_2966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2968 = 6'h2e == _myNewVec_19_T_3[5:0] ? myVec_46 : _GEN_2967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2969 = 6'h2f == _myNewVec_19_T_3[5:0] ? myVec_47 : _GEN_2968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2970 = 6'h30 == _myNewVec_19_T_3[5:0] ? myVec_48 : _GEN_2969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2971 = 6'h31 == _myNewVec_19_T_3[5:0] ? myVec_49 : _GEN_2970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2972 = 6'h32 == _myNewVec_19_T_3[5:0] ? myVec_50 : _GEN_2971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2973 = 6'h33 == _myNewVec_19_T_3[5:0] ? myVec_51 : _GEN_2972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2974 = 6'h34 == _myNewVec_19_T_3[5:0] ? myVec_52 : _GEN_2973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2975 = 6'h35 == _myNewVec_19_T_3[5:0] ? myVec_53 : _GEN_2974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2976 = 6'h36 == _myNewVec_19_T_3[5:0] ? myVec_54 : _GEN_2975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2977 = 6'h37 == _myNewVec_19_T_3[5:0] ? myVec_55 : _GEN_2976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2978 = 6'h38 == _myNewVec_19_T_3[5:0] ? myVec_56 : _GEN_2977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2979 = 6'h39 == _myNewVec_19_T_3[5:0] ? myVec_57 : _GEN_2978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2980 = 6'h3a == _myNewVec_19_T_3[5:0] ? myVec_58 : _GEN_2979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2981 = 6'h3b == _myNewVec_19_T_3[5:0] ? myVec_59 : _GEN_2980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2982 = 6'h3c == _myNewVec_19_T_3[5:0] ? myVec_60 : _GEN_2981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2983 = 6'h3d == _myNewVec_19_T_3[5:0] ? myVec_61 : _GEN_2982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2984 = 6'h3e == _myNewVec_19_T_3[5:0] ? myVec_62 : _GEN_2983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_19 = 6'h3f == _myNewVec_19_T_3[5:0] ? myVec_63 : _GEN_2984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_18_T_3 = _myNewVec_63_T_1 + 16'h2d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_2987 = 6'h1 == _myNewVec_18_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2988 = 6'h2 == _myNewVec_18_T_3[5:0] ? myVec_2 : _GEN_2987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2989 = 6'h3 == _myNewVec_18_T_3[5:0] ? myVec_3 : _GEN_2988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2990 = 6'h4 == _myNewVec_18_T_3[5:0] ? myVec_4 : _GEN_2989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2991 = 6'h5 == _myNewVec_18_T_3[5:0] ? myVec_5 : _GEN_2990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2992 = 6'h6 == _myNewVec_18_T_3[5:0] ? myVec_6 : _GEN_2991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2993 = 6'h7 == _myNewVec_18_T_3[5:0] ? myVec_7 : _GEN_2992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2994 = 6'h8 == _myNewVec_18_T_3[5:0] ? myVec_8 : _GEN_2993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2995 = 6'h9 == _myNewVec_18_T_3[5:0] ? myVec_9 : _GEN_2994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2996 = 6'ha == _myNewVec_18_T_3[5:0] ? myVec_10 : _GEN_2995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2997 = 6'hb == _myNewVec_18_T_3[5:0] ? myVec_11 : _GEN_2996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2998 = 6'hc == _myNewVec_18_T_3[5:0] ? myVec_12 : _GEN_2997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_2999 = 6'hd == _myNewVec_18_T_3[5:0] ? myVec_13 : _GEN_2998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3000 = 6'he == _myNewVec_18_T_3[5:0] ? myVec_14 : _GEN_2999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3001 = 6'hf == _myNewVec_18_T_3[5:0] ? myVec_15 : _GEN_3000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3002 = 6'h10 == _myNewVec_18_T_3[5:0] ? myVec_16 : _GEN_3001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3003 = 6'h11 == _myNewVec_18_T_3[5:0] ? myVec_17 : _GEN_3002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3004 = 6'h12 == _myNewVec_18_T_3[5:0] ? myVec_18 : _GEN_3003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3005 = 6'h13 == _myNewVec_18_T_3[5:0] ? myVec_19 : _GEN_3004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3006 = 6'h14 == _myNewVec_18_T_3[5:0] ? myVec_20 : _GEN_3005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3007 = 6'h15 == _myNewVec_18_T_3[5:0] ? myVec_21 : _GEN_3006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3008 = 6'h16 == _myNewVec_18_T_3[5:0] ? myVec_22 : _GEN_3007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3009 = 6'h17 == _myNewVec_18_T_3[5:0] ? myVec_23 : _GEN_3008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3010 = 6'h18 == _myNewVec_18_T_3[5:0] ? myVec_24 : _GEN_3009; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3011 = 6'h19 == _myNewVec_18_T_3[5:0] ? myVec_25 : _GEN_3010; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3012 = 6'h1a == _myNewVec_18_T_3[5:0] ? myVec_26 : _GEN_3011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3013 = 6'h1b == _myNewVec_18_T_3[5:0] ? myVec_27 : _GEN_3012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3014 = 6'h1c == _myNewVec_18_T_3[5:0] ? myVec_28 : _GEN_3013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3015 = 6'h1d == _myNewVec_18_T_3[5:0] ? myVec_29 : _GEN_3014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3016 = 6'h1e == _myNewVec_18_T_3[5:0] ? myVec_30 : _GEN_3015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3017 = 6'h1f == _myNewVec_18_T_3[5:0] ? myVec_31 : _GEN_3016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3018 = 6'h20 == _myNewVec_18_T_3[5:0] ? myVec_32 : _GEN_3017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3019 = 6'h21 == _myNewVec_18_T_3[5:0] ? myVec_33 : _GEN_3018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3020 = 6'h22 == _myNewVec_18_T_3[5:0] ? myVec_34 : _GEN_3019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3021 = 6'h23 == _myNewVec_18_T_3[5:0] ? myVec_35 : _GEN_3020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3022 = 6'h24 == _myNewVec_18_T_3[5:0] ? myVec_36 : _GEN_3021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3023 = 6'h25 == _myNewVec_18_T_3[5:0] ? myVec_37 : _GEN_3022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3024 = 6'h26 == _myNewVec_18_T_3[5:0] ? myVec_38 : _GEN_3023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3025 = 6'h27 == _myNewVec_18_T_3[5:0] ? myVec_39 : _GEN_3024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3026 = 6'h28 == _myNewVec_18_T_3[5:0] ? myVec_40 : _GEN_3025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3027 = 6'h29 == _myNewVec_18_T_3[5:0] ? myVec_41 : _GEN_3026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3028 = 6'h2a == _myNewVec_18_T_3[5:0] ? myVec_42 : _GEN_3027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3029 = 6'h2b == _myNewVec_18_T_3[5:0] ? myVec_43 : _GEN_3028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3030 = 6'h2c == _myNewVec_18_T_3[5:0] ? myVec_44 : _GEN_3029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3031 = 6'h2d == _myNewVec_18_T_3[5:0] ? myVec_45 : _GEN_3030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3032 = 6'h2e == _myNewVec_18_T_3[5:0] ? myVec_46 : _GEN_3031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3033 = 6'h2f == _myNewVec_18_T_3[5:0] ? myVec_47 : _GEN_3032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3034 = 6'h30 == _myNewVec_18_T_3[5:0] ? myVec_48 : _GEN_3033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3035 = 6'h31 == _myNewVec_18_T_3[5:0] ? myVec_49 : _GEN_3034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3036 = 6'h32 == _myNewVec_18_T_3[5:0] ? myVec_50 : _GEN_3035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3037 = 6'h33 == _myNewVec_18_T_3[5:0] ? myVec_51 : _GEN_3036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3038 = 6'h34 == _myNewVec_18_T_3[5:0] ? myVec_52 : _GEN_3037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3039 = 6'h35 == _myNewVec_18_T_3[5:0] ? myVec_53 : _GEN_3038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3040 = 6'h36 == _myNewVec_18_T_3[5:0] ? myVec_54 : _GEN_3039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3041 = 6'h37 == _myNewVec_18_T_3[5:0] ? myVec_55 : _GEN_3040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3042 = 6'h38 == _myNewVec_18_T_3[5:0] ? myVec_56 : _GEN_3041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3043 = 6'h39 == _myNewVec_18_T_3[5:0] ? myVec_57 : _GEN_3042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3044 = 6'h3a == _myNewVec_18_T_3[5:0] ? myVec_58 : _GEN_3043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3045 = 6'h3b == _myNewVec_18_T_3[5:0] ? myVec_59 : _GEN_3044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3046 = 6'h3c == _myNewVec_18_T_3[5:0] ? myVec_60 : _GEN_3045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3047 = 6'h3d == _myNewVec_18_T_3[5:0] ? myVec_61 : _GEN_3046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3048 = 6'h3e == _myNewVec_18_T_3[5:0] ? myVec_62 : _GEN_3047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_18 = 6'h3f == _myNewVec_18_T_3[5:0] ? myVec_63 : _GEN_3048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_17_T_3 = _myNewVec_63_T_1 + 16'h2e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3051 = 6'h1 == _myNewVec_17_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3052 = 6'h2 == _myNewVec_17_T_3[5:0] ? myVec_2 : _GEN_3051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3053 = 6'h3 == _myNewVec_17_T_3[5:0] ? myVec_3 : _GEN_3052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3054 = 6'h4 == _myNewVec_17_T_3[5:0] ? myVec_4 : _GEN_3053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3055 = 6'h5 == _myNewVec_17_T_3[5:0] ? myVec_5 : _GEN_3054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3056 = 6'h6 == _myNewVec_17_T_3[5:0] ? myVec_6 : _GEN_3055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3057 = 6'h7 == _myNewVec_17_T_3[5:0] ? myVec_7 : _GEN_3056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3058 = 6'h8 == _myNewVec_17_T_3[5:0] ? myVec_8 : _GEN_3057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3059 = 6'h9 == _myNewVec_17_T_3[5:0] ? myVec_9 : _GEN_3058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3060 = 6'ha == _myNewVec_17_T_3[5:0] ? myVec_10 : _GEN_3059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3061 = 6'hb == _myNewVec_17_T_3[5:0] ? myVec_11 : _GEN_3060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3062 = 6'hc == _myNewVec_17_T_3[5:0] ? myVec_12 : _GEN_3061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3063 = 6'hd == _myNewVec_17_T_3[5:0] ? myVec_13 : _GEN_3062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3064 = 6'he == _myNewVec_17_T_3[5:0] ? myVec_14 : _GEN_3063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3065 = 6'hf == _myNewVec_17_T_3[5:0] ? myVec_15 : _GEN_3064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3066 = 6'h10 == _myNewVec_17_T_3[5:0] ? myVec_16 : _GEN_3065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3067 = 6'h11 == _myNewVec_17_T_3[5:0] ? myVec_17 : _GEN_3066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3068 = 6'h12 == _myNewVec_17_T_3[5:0] ? myVec_18 : _GEN_3067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3069 = 6'h13 == _myNewVec_17_T_3[5:0] ? myVec_19 : _GEN_3068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3070 = 6'h14 == _myNewVec_17_T_3[5:0] ? myVec_20 : _GEN_3069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3071 = 6'h15 == _myNewVec_17_T_3[5:0] ? myVec_21 : _GEN_3070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3072 = 6'h16 == _myNewVec_17_T_3[5:0] ? myVec_22 : _GEN_3071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3073 = 6'h17 == _myNewVec_17_T_3[5:0] ? myVec_23 : _GEN_3072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3074 = 6'h18 == _myNewVec_17_T_3[5:0] ? myVec_24 : _GEN_3073; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3075 = 6'h19 == _myNewVec_17_T_3[5:0] ? myVec_25 : _GEN_3074; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3076 = 6'h1a == _myNewVec_17_T_3[5:0] ? myVec_26 : _GEN_3075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3077 = 6'h1b == _myNewVec_17_T_3[5:0] ? myVec_27 : _GEN_3076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3078 = 6'h1c == _myNewVec_17_T_3[5:0] ? myVec_28 : _GEN_3077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3079 = 6'h1d == _myNewVec_17_T_3[5:0] ? myVec_29 : _GEN_3078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3080 = 6'h1e == _myNewVec_17_T_3[5:0] ? myVec_30 : _GEN_3079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3081 = 6'h1f == _myNewVec_17_T_3[5:0] ? myVec_31 : _GEN_3080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3082 = 6'h20 == _myNewVec_17_T_3[5:0] ? myVec_32 : _GEN_3081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3083 = 6'h21 == _myNewVec_17_T_3[5:0] ? myVec_33 : _GEN_3082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3084 = 6'h22 == _myNewVec_17_T_3[5:0] ? myVec_34 : _GEN_3083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3085 = 6'h23 == _myNewVec_17_T_3[5:0] ? myVec_35 : _GEN_3084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3086 = 6'h24 == _myNewVec_17_T_3[5:0] ? myVec_36 : _GEN_3085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3087 = 6'h25 == _myNewVec_17_T_3[5:0] ? myVec_37 : _GEN_3086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3088 = 6'h26 == _myNewVec_17_T_3[5:0] ? myVec_38 : _GEN_3087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3089 = 6'h27 == _myNewVec_17_T_3[5:0] ? myVec_39 : _GEN_3088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3090 = 6'h28 == _myNewVec_17_T_3[5:0] ? myVec_40 : _GEN_3089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3091 = 6'h29 == _myNewVec_17_T_3[5:0] ? myVec_41 : _GEN_3090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3092 = 6'h2a == _myNewVec_17_T_3[5:0] ? myVec_42 : _GEN_3091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3093 = 6'h2b == _myNewVec_17_T_3[5:0] ? myVec_43 : _GEN_3092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3094 = 6'h2c == _myNewVec_17_T_3[5:0] ? myVec_44 : _GEN_3093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3095 = 6'h2d == _myNewVec_17_T_3[5:0] ? myVec_45 : _GEN_3094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3096 = 6'h2e == _myNewVec_17_T_3[5:0] ? myVec_46 : _GEN_3095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3097 = 6'h2f == _myNewVec_17_T_3[5:0] ? myVec_47 : _GEN_3096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3098 = 6'h30 == _myNewVec_17_T_3[5:0] ? myVec_48 : _GEN_3097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3099 = 6'h31 == _myNewVec_17_T_3[5:0] ? myVec_49 : _GEN_3098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3100 = 6'h32 == _myNewVec_17_T_3[5:0] ? myVec_50 : _GEN_3099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3101 = 6'h33 == _myNewVec_17_T_3[5:0] ? myVec_51 : _GEN_3100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3102 = 6'h34 == _myNewVec_17_T_3[5:0] ? myVec_52 : _GEN_3101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3103 = 6'h35 == _myNewVec_17_T_3[5:0] ? myVec_53 : _GEN_3102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3104 = 6'h36 == _myNewVec_17_T_3[5:0] ? myVec_54 : _GEN_3103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3105 = 6'h37 == _myNewVec_17_T_3[5:0] ? myVec_55 : _GEN_3104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3106 = 6'h38 == _myNewVec_17_T_3[5:0] ? myVec_56 : _GEN_3105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3107 = 6'h39 == _myNewVec_17_T_3[5:0] ? myVec_57 : _GEN_3106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3108 = 6'h3a == _myNewVec_17_T_3[5:0] ? myVec_58 : _GEN_3107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3109 = 6'h3b == _myNewVec_17_T_3[5:0] ? myVec_59 : _GEN_3108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3110 = 6'h3c == _myNewVec_17_T_3[5:0] ? myVec_60 : _GEN_3109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3111 = 6'h3d == _myNewVec_17_T_3[5:0] ? myVec_61 : _GEN_3110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3112 = 6'h3e == _myNewVec_17_T_3[5:0] ? myVec_62 : _GEN_3111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_17 = 6'h3f == _myNewVec_17_T_3[5:0] ? myVec_63 : _GEN_3112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_16_T_3 = _myNewVec_63_T_1 + 16'h2f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3115 = 6'h1 == _myNewVec_16_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3116 = 6'h2 == _myNewVec_16_T_3[5:0] ? myVec_2 : _GEN_3115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3117 = 6'h3 == _myNewVec_16_T_3[5:0] ? myVec_3 : _GEN_3116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3118 = 6'h4 == _myNewVec_16_T_3[5:0] ? myVec_4 : _GEN_3117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3119 = 6'h5 == _myNewVec_16_T_3[5:0] ? myVec_5 : _GEN_3118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3120 = 6'h6 == _myNewVec_16_T_3[5:0] ? myVec_6 : _GEN_3119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3121 = 6'h7 == _myNewVec_16_T_3[5:0] ? myVec_7 : _GEN_3120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3122 = 6'h8 == _myNewVec_16_T_3[5:0] ? myVec_8 : _GEN_3121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3123 = 6'h9 == _myNewVec_16_T_3[5:0] ? myVec_9 : _GEN_3122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3124 = 6'ha == _myNewVec_16_T_3[5:0] ? myVec_10 : _GEN_3123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3125 = 6'hb == _myNewVec_16_T_3[5:0] ? myVec_11 : _GEN_3124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3126 = 6'hc == _myNewVec_16_T_3[5:0] ? myVec_12 : _GEN_3125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3127 = 6'hd == _myNewVec_16_T_3[5:0] ? myVec_13 : _GEN_3126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3128 = 6'he == _myNewVec_16_T_3[5:0] ? myVec_14 : _GEN_3127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3129 = 6'hf == _myNewVec_16_T_3[5:0] ? myVec_15 : _GEN_3128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3130 = 6'h10 == _myNewVec_16_T_3[5:0] ? myVec_16 : _GEN_3129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3131 = 6'h11 == _myNewVec_16_T_3[5:0] ? myVec_17 : _GEN_3130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3132 = 6'h12 == _myNewVec_16_T_3[5:0] ? myVec_18 : _GEN_3131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3133 = 6'h13 == _myNewVec_16_T_3[5:0] ? myVec_19 : _GEN_3132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3134 = 6'h14 == _myNewVec_16_T_3[5:0] ? myVec_20 : _GEN_3133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3135 = 6'h15 == _myNewVec_16_T_3[5:0] ? myVec_21 : _GEN_3134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3136 = 6'h16 == _myNewVec_16_T_3[5:0] ? myVec_22 : _GEN_3135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3137 = 6'h17 == _myNewVec_16_T_3[5:0] ? myVec_23 : _GEN_3136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3138 = 6'h18 == _myNewVec_16_T_3[5:0] ? myVec_24 : _GEN_3137; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3139 = 6'h19 == _myNewVec_16_T_3[5:0] ? myVec_25 : _GEN_3138; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3140 = 6'h1a == _myNewVec_16_T_3[5:0] ? myVec_26 : _GEN_3139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3141 = 6'h1b == _myNewVec_16_T_3[5:0] ? myVec_27 : _GEN_3140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3142 = 6'h1c == _myNewVec_16_T_3[5:0] ? myVec_28 : _GEN_3141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3143 = 6'h1d == _myNewVec_16_T_3[5:0] ? myVec_29 : _GEN_3142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3144 = 6'h1e == _myNewVec_16_T_3[5:0] ? myVec_30 : _GEN_3143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3145 = 6'h1f == _myNewVec_16_T_3[5:0] ? myVec_31 : _GEN_3144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3146 = 6'h20 == _myNewVec_16_T_3[5:0] ? myVec_32 : _GEN_3145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3147 = 6'h21 == _myNewVec_16_T_3[5:0] ? myVec_33 : _GEN_3146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3148 = 6'h22 == _myNewVec_16_T_3[5:0] ? myVec_34 : _GEN_3147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3149 = 6'h23 == _myNewVec_16_T_3[5:0] ? myVec_35 : _GEN_3148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3150 = 6'h24 == _myNewVec_16_T_3[5:0] ? myVec_36 : _GEN_3149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3151 = 6'h25 == _myNewVec_16_T_3[5:0] ? myVec_37 : _GEN_3150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3152 = 6'h26 == _myNewVec_16_T_3[5:0] ? myVec_38 : _GEN_3151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3153 = 6'h27 == _myNewVec_16_T_3[5:0] ? myVec_39 : _GEN_3152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3154 = 6'h28 == _myNewVec_16_T_3[5:0] ? myVec_40 : _GEN_3153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3155 = 6'h29 == _myNewVec_16_T_3[5:0] ? myVec_41 : _GEN_3154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3156 = 6'h2a == _myNewVec_16_T_3[5:0] ? myVec_42 : _GEN_3155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3157 = 6'h2b == _myNewVec_16_T_3[5:0] ? myVec_43 : _GEN_3156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3158 = 6'h2c == _myNewVec_16_T_3[5:0] ? myVec_44 : _GEN_3157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3159 = 6'h2d == _myNewVec_16_T_3[5:0] ? myVec_45 : _GEN_3158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3160 = 6'h2e == _myNewVec_16_T_3[5:0] ? myVec_46 : _GEN_3159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3161 = 6'h2f == _myNewVec_16_T_3[5:0] ? myVec_47 : _GEN_3160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3162 = 6'h30 == _myNewVec_16_T_3[5:0] ? myVec_48 : _GEN_3161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3163 = 6'h31 == _myNewVec_16_T_3[5:0] ? myVec_49 : _GEN_3162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3164 = 6'h32 == _myNewVec_16_T_3[5:0] ? myVec_50 : _GEN_3163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3165 = 6'h33 == _myNewVec_16_T_3[5:0] ? myVec_51 : _GEN_3164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3166 = 6'h34 == _myNewVec_16_T_3[5:0] ? myVec_52 : _GEN_3165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3167 = 6'h35 == _myNewVec_16_T_3[5:0] ? myVec_53 : _GEN_3166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3168 = 6'h36 == _myNewVec_16_T_3[5:0] ? myVec_54 : _GEN_3167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3169 = 6'h37 == _myNewVec_16_T_3[5:0] ? myVec_55 : _GEN_3168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3170 = 6'h38 == _myNewVec_16_T_3[5:0] ? myVec_56 : _GEN_3169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3171 = 6'h39 == _myNewVec_16_T_3[5:0] ? myVec_57 : _GEN_3170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3172 = 6'h3a == _myNewVec_16_T_3[5:0] ? myVec_58 : _GEN_3171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3173 = 6'h3b == _myNewVec_16_T_3[5:0] ? myVec_59 : _GEN_3172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3174 = 6'h3c == _myNewVec_16_T_3[5:0] ? myVec_60 : _GEN_3173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3175 = 6'h3d == _myNewVec_16_T_3[5:0] ? myVec_61 : _GEN_3174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3176 = 6'h3e == _myNewVec_16_T_3[5:0] ? myVec_62 : _GEN_3175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_16 = 6'h3f == _myNewVec_16_T_3[5:0] ? myVec_63 : _GEN_3176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_hi_lo = {myNewVec_23,myNewVec_22,myNewVec_21,myNewVec_20,myNewVec_19,myNewVec_18,myNewVec_17
    ,myNewVec_16}; // @[hh_datapath_chisel.scala 238:27]
  wire [15:0] _myNewVec_15_T_3 = _myNewVec_63_T_1 + 16'h30; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3179 = 6'h1 == _myNewVec_15_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3180 = 6'h2 == _myNewVec_15_T_3[5:0] ? myVec_2 : _GEN_3179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3181 = 6'h3 == _myNewVec_15_T_3[5:0] ? myVec_3 : _GEN_3180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3182 = 6'h4 == _myNewVec_15_T_3[5:0] ? myVec_4 : _GEN_3181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3183 = 6'h5 == _myNewVec_15_T_3[5:0] ? myVec_5 : _GEN_3182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3184 = 6'h6 == _myNewVec_15_T_3[5:0] ? myVec_6 : _GEN_3183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3185 = 6'h7 == _myNewVec_15_T_3[5:0] ? myVec_7 : _GEN_3184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3186 = 6'h8 == _myNewVec_15_T_3[5:0] ? myVec_8 : _GEN_3185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3187 = 6'h9 == _myNewVec_15_T_3[5:0] ? myVec_9 : _GEN_3186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3188 = 6'ha == _myNewVec_15_T_3[5:0] ? myVec_10 : _GEN_3187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3189 = 6'hb == _myNewVec_15_T_3[5:0] ? myVec_11 : _GEN_3188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3190 = 6'hc == _myNewVec_15_T_3[5:0] ? myVec_12 : _GEN_3189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3191 = 6'hd == _myNewVec_15_T_3[5:0] ? myVec_13 : _GEN_3190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3192 = 6'he == _myNewVec_15_T_3[5:0] ? myVec_14 : _GEN_3191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3193 = 6'hf == _myNewVec_15_T_3[5:0] ? myVec_15 : _GEN_3192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3194 = 6'h10 == _myNewVec_15_T_3[5:0] ? myVec_16 : _GEN_3193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3195 = 6'h11 == _myNewVec_15_T_3[5:0] ? myVec_17 : _GEN_3194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3196 = 6'h12 == _myNewVec_15_T_3[5:0] ? myVec_18 : _GEN_3195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3197 = 6'h13 == _myNewVec_15_T_3[5:0] ? myVec_19 : _GEN_3196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3198 = 6'h14 == _myNewVec_15_T_3[5:0] ? myVec_20 : _GEN_3197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3199 = 6'h15 == _myNewVec_15_T_3[5:0] ? myVec_21 : _GEN_3198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3200 = 6'h16 == _myNewVec_15_T_3[5:0] ? myVec_22 : _GEN_3199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3201 = 6'h17 == _myNewVec_15_T_3[5:0] ? myVec_23 : _GEN_3200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3202 = 6'h18 == _myNewVec_15_T_3[5:0] ? myVec_24 : _GEN_3201; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3203 = 6'h19 == _myNewVec_15_T_3[5:0] ? myVec_25 : _GEN_3202; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3204 = 6'h1a == _myNewVec_15_T_3[5:0] ? myVec_26 : _GEN_3203; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3205 = 6'h1b == _myNewVec_15_T_3[5:0] ? myVec_27 : _GEN_3204; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3206 = 6'h1c == _myNewVec_15_T_3[5:0] ? myVec_28 : _GEN_3205; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3207 = 6'h1d == _myNewVec_15_T_3[5:0] ? myVec_29 : _GEN_3206; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3208 = 6'h1e == _myNewVec_15_T_3[5:0] ? myVec_30 : _GEN_3207; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3209 = 6'h1f == _myNewVec_15_T_3[5:0] ? myVec_31 : _GEN_3208; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3210 = 6'h20 == _myNewVec_15_T_3[5:0] ? myVec_32 : _GEN_3209; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3211 = 6'h21 == _myNewVec_15_T_3[5:0] ? myVec_33 : _GEN_3210; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3212 = 6'h22 == _myNewVec_15_T_3[5:0] ? myVec_34 : _GEN_3211; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3213 = 6'h23 == _myNewVec_15_T_3[5:0] ? myVec_35 : _GEN_3212; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3214 = 6'h24 == _myNewVec_15_T_3[5:0] ? myVec_36 : _GEN_3213; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3215 = 6'h25 == _myNewVec_15_T_3[5:0] ? myVec_37 : _GEN_3214; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3216 = 6'h26 == _myNewVec_15_T_3[5:0] ? myVec_38 : _GEN_3215; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3217 = 6'h27 == _myNewVec_15_T_3[5:0] ? myVec_39 : _GEN_3216; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3218 = 6'h28 == _myNewVec_15_T_3[5:0] ? myVec_40 : _GEN_3217; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3219 = 6'h29 == _myNewVec_15_T_3[5:0] ? myVec_41 : _GEN_3218; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3220 = 6'h2a == _myNewVec_15_T_3[5:0] ? myVec_42 : _GEN_3219; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3221 = 6'h2b == _myNewVec_15_T_3[5:0] ? myVec_43 : _GEN_3220; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3222 = 6'h2c == _myNewVec_15_T_3[5:0] ? myVec_44 : _GEN_3221; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3223 = 6'h2d == _myNewVec_15_T_3[5:0] ? myVec_45 : _GEN_3222; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3224 = 6'h2e == _myNewVec_15_T_3[5:0] ? myVec_46 : _GEN_3223; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3225 = 6'h2f == _myNewVec_15_T_3[5:0] ? myVec_47 : _GEN_3224; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3226 = 6'h30 == _myNewVec_15_T_3[5:0] ? myVec_48 : _GEN_3225; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3227 = 6'h31 == _myNewVec_15_T_3[5:0] ? myVec_49 : _GEN_3226; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3228 = 6'h32 == _myNewVec_15_T_3[5:0] ? myVec_50 : _GEN_3227; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3229 = 6'h33 == _myNewVec_15_T_3[5:0] ? myVec_51 : _GEN_3228; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3230 = 6'h34 == _myNewVec_15_T_3[5:0] ? myVec_52 : _GEN_3229; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3231 = 6'h35 == _myNewVec_15_T_3[5:0] ? myVec_53 : _GEN_3230; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3232 = 6'h36 == _myNewVec_15_T_3[5:0] ? myVec_54 : _GEN_3231; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3233 = 6'h37 == _myNewVec_15_T_3[5:0] ? myVec_55 : _GEN_3232; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3234 = 6'h38 == _myNewVec_15_T_3[5:0] ? myVec_56 : _GEN_3233; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3235 = 6'h39 == _myNewVec_15_T_3[5:0] ? myVec_57 : _GEN_3234; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3236 = 6'h3a == _myNewVec_15_T_3[5:0] ? myVec_58 : _GEN_3235; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3237 = 6'h3b == _myNewVec_15_T_3[5:0] ? myVec_59 : _GEN_3236; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3238 = 6'h3c == _myNewVec_15_T_3[5:0] ? myVec_60 : _GEN_3237; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3239 = 6'h3d == _myNewVec_15_T_3[5:0] ? myVec_61 : _GEN_3238; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3240 = 6'h3e == _myNewVec_15_T_3[5:0] ? myVec_62 : _GEN_3239; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_15 = 6'h3f == _myNewVec_15_T_3[5:0] ? myVec_63 : _GEN_3240; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_14_T_3 = _myNewVec_63_T_1 + 16'h31; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3243 = 6'h1 == _myNewVec_14_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3244 = 6'h2 == _myNewVec_14_T_3[5:0] ? myVec_2 : _GEN_3243; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3245 = 6'h3 == _myNewVec_14_T_3[5:0] ? myVec_3 : _GEN_3244; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3246 = 6'h4 == _myNewVec_14_T_3[5:0] ? myVec_4 : _GEN_3245; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3247 = 6'h5 == _myNewVec_14_T_3[5:0] ? myVec_5 : _GEN_3246; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3248 = 6'h6 == _myNewVec_14_T_3[5:0] ? myVec_6 : _GEN_3247; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3249 = 6'h7 == _myNewVec_14_T_3[5:0] ? myVec_7 : _GEN_3248; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3250 = 6'h8 == _myNewVec_14_T_3[5:0] ? myVec_8 : _GEN_3249; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3251 = 6'h9 == _myNewVec_14_T_3[5:0] ? myVec_9 : _GEN_3250; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3252 = 6'ha == _myNewVec_14_T_3[5:0] ? myVec_10 : _GEN_3251; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3253 = 6'hb == _myNewVec_14_T_3[5:0] ? myVec_11 : _GEN_3252; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3254 = 6'hc == _myNewVec_14_T_3[5:0] ? myVec_12 : _GEN_3253; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3255 = 6'hd == _myNewVec_14_T_3[5:0] ? myVec_13 : _GEN_3254; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3256 = 6'he == _myNewVec_14_T_3[5:0] ? myVec_14 : _GEN_3255; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3257 = 6'hf == _myNewVec_14_T_3[5:0] ? myVec_15 : _GEN_3256; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3258 = 6'h10 == _myNewVec_14_T_3[5:0] ? myVec_16 : _GEN_3257; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3259 = 6'h11 == _myNewVec_14_T_3[5:0] ? myVec_17 : _GEN_3258; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3260 = 6'h12 == _myNewVec_14_T_3[5:0] ? myVec_18 : _GEN_3259; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3261 = 6'h13 == _myNewVec_14_T_3[5:0] ? myVec_19 : _GEN_3260; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3262 = 6'h14 == _myNewVec_14_T_3[5:0] ? myVec_20 : _GEN_3261; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3263 = 6'h15 == _myNewVec_14_T_3[5:0] ? myVec_21 : _GEN_3262; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3264 = 6'h16 == _myNewVec_14_T_3[5:0] ? myVec_22 : _GEN_3263; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3265 = 6'h17 == _myNewVec_14_T_3[5:0] ? myVec_23 : _GEN_3264; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3266 = 6'h18 == _myNewVec_14_T_3[5:0] ? myVec_24 : _GEN_3265; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3267 = 6'h19 == _myNewVec_14_T_3[5:0] ? myVec_25 : _GEN_3266; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3268 = 6'h1a == _myNewVec_14_T_3[5:0] ? myVec_26 : _GEN_3267; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3269 = 6'h1b == _myNewVec_14_T_3[5:0] ? myVec_27 : _GEN_3268; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3270 = 6'h1c == _myNewVec_14_T_3[5:0] ? myVec_28 : _GEN_3269; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3271 = 6'h1d == _myNewVec_14_T_3[5:0] ? myVec_29 : _GEN_3270; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3272 = 6'h1e == _myNewVec_14_T_3[5:0] ? myVec_30 : _GEN_3271; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3273 = 6'h1f == _myNewVec_14_T_3[5:0] ? myVec_31 : _GEN_3272; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3274 = 6'h20 == _myNewVec_14_T_3[5:0] ? myVec_32 : _GEN_3273; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3275 = 6'h21 == _myNewVec_14_T_3[5:0] ? myVec_33 : _GEN_3274; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3276 = 6'h22 == _myNewVec_14_T_3[5:0] ? myVec_34 : _GEN_3275; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3277 = 6'h23 == _myNewVec_14_T_3[5:0] ? myVec_35 : _GEN_3276; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3278 = 6'h24 == _myNewVec_14_T_3[5:0] ? myVec_36 : _GEN_3277; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3279 = 6'h25 == _myNewVec_14_T_3[5:0] ? myVec_37 : _GEN_3278; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3280 = 6'h26 == _myNewVec_14_T_3[5:0] ? myVec_38 : _GEN_3279; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3281 = 6'h27 == _myNewVec_14_T_3[5:0] ? myVec_39 : _GEN_3280; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3282 = 6'h28 == _myNewVec_14_T_3[5:0] ? myVec_40 : _GEN_3281; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3283 = 6'h29 == _myNewVec_14_T_3[5:0] ? myVec_41 : _GEN_3282; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3284 = 6'h2a == _myNewVec_14_T_3[5:0] ? myVec_42 : _GEN_3283; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3285 = 6'h2b == _myNewVec_14_T_3[5:0] ? myVec_43 : _GEN_3284; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3286 = 6'h2c == _myNewVec_14_T_3[5:0] ? myVec_44 : _GEN_3285; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3287 = 6'h2d == _myNewVec_14_T_3[5:0] ? myVec_45 : _GEN_3286; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3288 = 6'h2e == _myNewVec_14_T_3[5:0] ? myVec_46 : _GEN_3287; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3289 = 6'h2f == _myNewVec_14_T_3[5:0] ? myVec_47 : _GEN_3288; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3290 = 6'h30 == _myNewVec_14_T_3[5:0] ? myVec_48 : _GEN_3289; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3291 = 6'h31 == _myNewVec_14_T_3[5:0] ? myVec_49 : _GEN_3290; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3292 = 6'h32 == _myNewVec_14_T_3[5:0] ? myVec_50 : _GEN_3291; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3293 = 6'h33 == _myNewVec_14_T_3[5:0] ? myVec_51 : _GEN_3292; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3294 = 6'h34 == _myNewVec_14_T_3[5:0] ? myVec_52 : _GEN_3293; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3295 = 6'h35 == _myNewVec_14_T_3[5:0] ? myVec_53 : _GEN_3294; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3296 = 6'h36 == _myNewVec_14_T_3[5:0] ? myVec_54 : _GEN_3295; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3297 = 6'h37 == _myNewVec_14_T_3[5:0] ? myVec_55 : _GEN_3296; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3298 = 6'h38 == _myNewVec_14_T_3[5:0] ? myVec_56 : _GEN_3297; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3299 = 6'h39 == _myNewVec_14_T_3[5:0] ? myVec_57 : _GEN_3298; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3300 = 6'h3a == _myNewVec_14_T_3[5:0] ? myVec_58 : _GEN_3299; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3301 = 6'h3b == _myNewVec_14_T_3[5:0] ? myVec_59 : _GEN_3300; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3302 = 6'h3c == _myNewVec_14_T_3[5:0] ? myVec_60 : _GEN_3301; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3303 = 6'h3d == _myNewVec_14_T_3[5:0] ? myVec_61 : _GEN_3302; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3304 = 6'h3e == _myNewVec_14_T_3[5:0] ? myVec_62 : _GEN_3303; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_14 = 6'h3f == _myNewVec_14_T_3[5:0] ? myVec_63 : _GEN_3304; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_13_T_3 = _myNewVec_63_T_1 + 16'h32; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3307 = 6'h1 == _myNewVec_13_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3308 = 6'h2 == _myNewVec_13_T_3[5:0] ? myVec_2 : _GEN_3307; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3309 = 6'h3 == _myNewVec_13_T_3[5:0] ? myVec_3 : _GEN_3308; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3310 = 6'h4 == _myNewVec_13_T_3[5:0] ? myVec_4 : _GEN_3309; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3311 = 6'h5 == _myNewVec_13_T_3[5:0] ? myVec_5 : _GEN_3310; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3312 = 6'h6 == _myNewVec_13_T_3[5:0] ? myVec_6 : _GEN_3311; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3313 = 6'h7 == _myNewVec_13_T_3[5:0] ? myVec_7 : _GEN_3312; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3314 = 6'h8 == _myNewVec_13_T_3[5:0] ? myVec_8 : _GEN_3313; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3315 = 6'h9 == _myNewVec_13_T_3[5:0] ? myVec_9 : _GEN_3314; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3316 = 6'ha == _myNewVec_13_T_3[5:0] ? myVec_10 : _GEN_3315; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3317 = 6'hb == _myNewVec_13_T_3[5:0] ? myVec_11 : _GEN_3316; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3318 = 6'hc == _myNewVec_13_T_3[5:0] ? myVec_12 : _GEN_3317; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3319 = 6'hd == _myNewVec_13_T_3[5:0] ? myVec_13 : _GEN_3318; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3320 = 6'he == _myNewVec_13_T_3[5:0] ? myVec_14 : _GEN_3319; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3321 = 6'hf == _myNewVec_13_T_3[5:0] ? myVec_15 : _GEN_3320; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3322 = 6'h10 == _myNewVec_13_T_3[5:0] ? myVec_16 : _GEN_3321; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3323 = 6'h11 == _myNewVec_13_T_3[5:0] ? myVec_17 : _GEN_3322; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3324 = 6'h12 == _myNewVec_13_T_3[5:0] ? myVec_18 : _GEN_3323; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3325 = 6'h13 == _myNewVec_13_T_3[5:0] ? myVec_19 : _GEN_3324; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3326 = 6'h14 == _myNewVec_13_T_3[5:0] ? myVec_20 : _GEN_3325; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3327 = 6'h15 == _myNewVec_13_T_3[5:0] ? myVec_21 : _GEN_3326; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3328 = 6'h16 == _myNewVec_13_T_3[5:0] ? myVec_22 : _GEN_3327; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3329 = 6'h17 == _myNewVec_13_T_3[5:0] ? myVec_23 : _GEN_3328; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3330 = 6'h18 == _myNewVec_13_T_3[5:0] ? myVec_24 : _GEN_3329; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3331 = 6'h19 == _myNewVec_13_T_3[5:0] ? myVec_25 : _GEN_3330; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3332 = 6'h1a == _myNewVec_13_T_3[5:0] ? myVec_26 : _GEN_3331; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3333 = 6'h1b == _myNewVec_13_T_3[5:0] ? myVec_27 : _GEN_3332; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3334 = 6'h1c == _myNewVec_13_T_3[5:0] ? myVec_28 : _GEN_3333; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3335 = 6'h1d == _myNewVec_13_T_3[5:0] ? myVec_29 : _GEN_3334; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3336 = 6'h1e == _myNewVec_13_T_3[5:0] ? myVec_30 : _GEN_3335; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3337 = 6'h1f == _myNewVec_13_T_3[5:0] ? myVec_31 : _GEN_3336; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3338 = 6'h20 == _myNewVec_13_T_3[5:0] ? myVec_32 : _GEN_3337; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3339 = 6'h21 == _myNewVec_13_T_3[5:0] ? myVec_33 : _GEN_3338; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3340 = 6'h22 == _myNewVec_13_T_3[5:0] ? myVec_34 : _GEN_3339; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3341 = 6'h23 == _myNewVec_13_T_3[5:0] ? myVec_35 : _GEN_3340; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3342 = 6'h24 == _myNewVec_13_T_3[5:0] ? myVec_36 : _GEN_3341; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3343 = 6'h25 == _myNewVec_13_T_3[5:0] ? myVec_37 : _GEN_3342; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3344 = 6'h26 == _myNewVec_13_T_3[5:0] ? myVec_38 : _GEN_3343; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3345 = 6'h27 == _myNewVec_13_T_3[5:0] ? myVec_39 : _GEN_3344; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3346 = 6'h28 == _myNewVec_13_T_3[5:0] ? myVec_40 : _GEN_3345; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3347 = 6'h29 == _myNewVec_13_T_3[5:0] ? myVec_41 : _GEN_3346; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3348 = 6'h2a == _myNewVec_13_T_3[5:0] ? myVec_42 : _GEN_3347; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3349 = 6'h2b == _myNewVec_13_T_3[5:0] ? myVec_43 : _GEN_3348; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3350 = 6'h2c == _myNewVec_13_T_3[5:0] ? myVec_44 : _GEN_3349; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3351 = 6'h2d == _myNewVec_13_T_3[5:0] ? myVec_45 : _GEN_3350; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3352 = 6'h2e == _myNewVec_13_T_3[5:0] ? myVec_46 : _GEN_3351; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3353 = 6'h2f == _myNewVec_13_T_3[5:0] ? myVec_47 : _GEN_3352; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3354 = 6'h30 == _myNewVec_13_T_3[5:0] ? myVec_48 : _GEN_3353; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3355 = 6'h31 == _myNewVec_13_T_3[5:0] ? myVec_49 : _GEN_3354; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3356 = 6'h32 == _myNewVec_13_T_3[5:0] ? myVec_50 : _GEN_3355; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3357 = 6'h33 == _myNewVec_13_T_3[5:0] ? myVec_51 : _GEN_3356; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3358 = 6'h34 == _myNewVec_13_T_3[5:0] ? myVec_52 : _GEN_3357; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3359 = 6'h35 == _myNewVec_13_T_3[5:0] ? myVec_53 : _GEN_3358; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3360 = 6'h36 == _myNewVec_13_T_3[5:0] ? myVec_54 : _GEN_3359; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3361 = 6'h37 == _myNewVec_13_T_3[5:0] ? myVec_55 : _GEN_3360; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3362 = 6'h38 == _myNewVec_13_T_3[5:0] ? myVec_56 : _GEN_3361; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3363 = 6'h39 == _myNewVec_13_T_3[5:0] ? myVec_57 : _GEN_3362; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3364 = 6'h3a == _myNewVec_13_T_3[5:0] ? myVec_58 : _GEN_3363; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3365 = 6'h3b == _myNewVec_13_T_3[5:0] ? myVec_59 : _GEN_3364; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3366 = 6'h3c == _myNewVec_13_T_3[5:0] ? myVec_60 : _GEN_3365; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3367 = 6'h3d == _myNewVec_13_T_3[5:0] ? myVec_61 : _GEN_3366; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3368 = 6'h3e == _myNewVec_13_T_3[5:0] ? myVec_62 : _GEN_3367; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_13 = 6'h3f == _myNewVec_13_T_3[5:0] ? myVec_63 : _GEN_3368; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_12_T_3 = _myNewVec_63_T_1 + 16'h33; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3371 = 6'h1 == _myNewVec_12_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3372 = 6'h2 == _myNewVec_12_T_3[5:0] ? myVec_2 : _GEN_3371; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3373 = 6'h3 == _myNewVec_12_T_3[5:0] ? myVec_3 : _GEN_3372; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3374 = 6'h4 == _myNewVec_12_T_3[5:0] ? myVec_4 : _GEN_3373; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3375 = 6'h5 == _myNewVec_12_T_3[5:0] ? myVec_5 : _GEN_3374; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3376 = 6'h6 == _myNewVec_12_T_3[5:0] ? myVec_6 : _GEN_3375; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3377 = 6'h7 == _myNewVec_12_T_3[5:0] ? myVec_7 : _GEN_3376; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3378 = 6'h8 == _myNewVec_12_T_3[5:0] ? myVec_8 : _GEN_3377; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3379 = 6'h9 == _myNewVec_12_T_3[5:0] ? myVec_9 : _GEN_3378; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3380 = 6'ha == _myNewVec_12_T_3[5:0] ? myVec_10 : _GEN_3379; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3381 = 6'hb == _myNewVec_12_T_3[5:0] ? myVec_11 : _GEN_3380; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3382 = 6'hc == _myNewVec_12_T_3[5:0] ? myVec_12 : _GEN_3381; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3383 = 6'hd == _myNewVec_12_T_3[5:0] ? myVec_13 : _GEN_3382; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3384 = 6'he == _myNewVec_12_T_3[5:0] ? myVec_14 : _GEN_3383; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3385 = 6'hf == _myNewVec_12_T_3[5:0] ? myVec_15 : _GEN_3384; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3386 = 6'h10 == _myNewVec_12_T_3[5:0] ? myVec_16 : _GEN_3385; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3387 = 6'h11 == _myNewVec_12_T_3[5:0] ? myVec_17 : _GEN_3386; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3388 = 6'h12 == _myNewVec_12_T_3[5:0] ? myVec_18 : _GEN_3387; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3389 = 6'h13 == _myNewVec_12_T_3[5:0] ? myVec_19 : _GEN_3388; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3390 = 6'h14 == _myNewVec_12_T_3[5:0] ? myVec_20 : _GEN_3389; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3391 = 6'h15 == _myNewVec_12_T_3[5:0] ? myVec_21 : _GEN_3390; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3392 = 6'h16 == _myNewVec_12_T_3[5:0] ? myVec_22 : _GEN_3391; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3393 = 6'h17 == _myNewVec_12_T_3[5:0] ? myVec_23 : _GEN_3392; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3394 = 6'h18 == _myNewVec_12_T_3[5:0] ? myVec_24 : _GEN_3393; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3395 = 6'h19 == _myNewVec_12_T_3[5:0] ? myVec_25 : _GEN_3394; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3396 = 6'h1a == _myNewVec_12_T_3[5:0] ? myVec_26 : _GEN_3395; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3397 = 6'h1b == _myNewVec_12_T_3[5:0] ? myVec_27 : _GEN_3396; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3398 = 6'h1c == _myNewVec_12_T_3[5:0] ? myVec_28 : _GEN_3397; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3399 = 6'h1d == _myNewVec_12_T_3[5:0] ? myVec_29 : _GEN_3398; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3400 = 6'h1e == _myNewVec_12_T_3[5:0] ? myVec_30 : _GEN_3399; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3401 = 6'h1f == _myNewVec_12_T_3[5:0] ? myVec_31 : _GEN_3400; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3402 = 6'h20 == _myNewVec_12_T_3[5:0] ? myVec_32 : _GEN_3401; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3403 = 6'h21 == _myNewVec_12_T_3[5:0] ? myVec_33 : _GEN_3402; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3404 = 6'h22 == _myNewVec_12_T_3[5:0] ? myVec_34 : _GEN_3403; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3405 = 6'h23 == _myNewVec_12_T_3[5:0] ? myVec_35 : _GEN_3404; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3406 = 6'h24 == _myNewVec_12_T_3[5:0] ? myVec_36 : _GEN_3405; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3407 = 6'h25 == _myNewVec_12_T_3[5:0] ? myVec_37 : _GEN_3406; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3408 = 6'h26 == _myNewVec_12_T_3[5:0] ? myVec_38 : _GEN_3407; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3409 = 6'h27 == _myNewVec_12_T_3[5:0] ? myVec_39 : _GEN_3408; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3410 = 6'h28 == _myNewVec_12_T_3[5:0] ? myVec_40 : _GEN_3409; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3411 = 6'h29 == _myNewVec_12_T_3[5:0] ? myVec_41 : _GEN_3410; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3412 = 6'h2a == _myNewVec_12_T_3[5:0] ? myVec_42 : _GEN_3411; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3413 = 6'h2b == _myNewVec_12_T_3[5:0] ? myVec_43 : _GEN_3412; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3414 = 6'h2c == _myNewVec_12_T_3[5:0] ? myVec_44 : _GEN_3413; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3415 = 6'h2d == _myNewVec_12_T_3[5:0] ? myVec_45 : _GEN_3414; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3416 = 6'h2e == _myNewVec_12_T_3[5:0] ? myVec_46 : _GEN_3415; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3417 = 6'h2f == _myNewVec_12_T_3[5:0] ? myVec_47 : _GEN_3416; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3418 = 6'h30 == _myNewVec_12_T_3[5:0] ? myVec_48 : _GEN_3417; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3419 = 6'h31 == _myNewVec_12_T_3[5:0] ? myVec_49 : _GEN_3418; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3420 = 6'h32 == _myNewVec_12_T_3[5:0] ? myVec_50 : _GEN_3419; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3421 = 6'h33 == _myNewVec_12_T_3[5:0] ? myVec_51 : _GEN_3420; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3422 = 6'h34 == _myNewVec_12_T_3[5:0] ? myVec_52 : _GEN_3421; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3423 = 6'h35 == _myNewVec_12_T_3[5:0] ? myVec_53 : _GEN_3422; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3424 = 6'h36 == _myNewVec_12_T_3[5:0] ? myVec_54 : _GEN_3423; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3425 = 6'h37 == _myNewVec_12_T_3[5:0] ? myVec_55 : _GEN_3424; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3426 = 6'h38 == _myNewVec_12_T_3[5:0] ? myVec_56 : _GEN_3425; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3427 = 6'h39 == _myNewVec_12_T_3[5:0] ? myVec_57 : _GEN_3426; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3428 = 6'h3a == _myNewVec_12_T_3[5:0] ? myVec_58 : _GEN_3427; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3429 = 6'h3b == _myNewVec_12_T_3[5:0] ? myVec_59 : _GEN_3428; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3430 = 6'h3c == _myNewVec_12_T_3[5:0] ? myVec_60 : _GEN_3429; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3431 = 6'h3d == _myNewVec_12_T_3[5:0] ? myVec_61 : _GEN_3430; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3432 = 6'h3e == _myNewVec_12_T_3[5:0] ? myVec_62 : _GEN_3431; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_12 = 6'h3f == _myNewVec_12_T_3[5:0] ? myVec_63 : _GEN_3432; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_11_T_3 = _myNewVec_63_T_1 + 16'h34; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3435 = 6'h1 == _myNewVec_11_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3436 = 6'h2 == _myNewVec_11_T_3[5:0] ? myVec_2 : _GEN_3435; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3437 = 6'h3 == _myNewVec_11_T_3[5:0] ? myVec_3 : _GEN_3436; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3438 = 6'h4 == _myNewVec_11_T_3[5:0] ? myVec_4 : _GEN_3437; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3439 = 6'h5 == _myNewVec_11_T_3[5:0] ? myVec_5 : _GEN_3438; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3440 = 6'h6 == _myNewVec_11_T_3[5:0] ? myVec_6 : _GEN_3439; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3441 = 6'h7 == _myNewVec_11_T_3[5:0] ? myVec_7 : _GEN_3440; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3442 = 6'h8 == _myNewVec_11_T_3[5:0] ? myVec_8 : _GEN_3441; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3443 = 6'h9 == _myNewVec_11_T_3[5:0] ? myVec_9 : _GEN_3442; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3444 = 6'ha == _myNewVec_11_T_3[5:0] ? myVec_10 : _GEN_3443; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3445 = 6'hb == _myNewVec_11_T_3[5:0] ? myVec_11 : _GEN_3444; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3446 = 6'hc == _myNewVec_11_T_3[5:0] ? myVec_12 : _GEN_3445; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3447 = 6'hd == _myNewVec_11_T_3[5:0] ? myVec_13 : _GEN_3446; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3448 = 6'he == _myNewVec_11_T_3[5:0] ? myVec_14 : _GEN_3447; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3449 = 6'hf == _myNewVec_11_T_3[5:0] ? myVec_15 : _GEN_3448; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3450 = 6'h10 == _myNewVec_11_T_3[5:0] ? myVec_16 : _GEN_3449; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3451 = 6'h11 == _myNewVec_11_T_3[5:0] ? myVec_17 : _GEN_3450; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3452 = 6'h12 == _myNewVec_11_T_3[5:0] ? myVec_18 : _GEN_3451; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3453 = 6'h13 == _myNewVec_11_T_3[5:0] ? myVec_19 : _GEN_3452; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3454 = 6'h14 == _myNewVec_11_T_3[5:0] ? myVec_20 : _GEN_3453; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3455 = 6'h15 == _myNewVec_11_T_3[5:0] ? myVec_21 : _GEN_3454; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3456 = 6'h16 == _myNewVec_11_T_3[5:0] ? myVec_22 : _GEN_3455; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3457 = 6'h17 == _myNewVec_11_T_3[5:0] ? myVec_23 : _GEN_3456; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3458 = 6'h18 == _myNewVec_11_T_3[5:0] ? myVec_24 : _GEN_3457; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3459 = 6'h19 == _myNewVec_11_T_3[5:0] ? myVec_25 : _GEN_3458; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3460 = 6'h1a == _myNewVec_11_T_3[5:0] ? myVec_26 : _GEN_3459; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3461 = 6'h1b == _myNewVec_11_T_3[5:0] ? myVec_27 : _GEN_3460; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3462 = 6'h1c == _myNewVec_11_T_3[5:0] ? myVec_28 : _GEN_3461; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3463 = 6'h1d == _myNewVec_11_T_3[5:0] ? myVec_29 : _GEN_3462; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3464 = 6'h1e == _myNewVec_11_T_3[5:0] ? myVec_30 : _GEN_3463; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3465 = 6'h1f == _myNewVec_11_T_3[5:0] ? myVec_31 : _GEN_3464; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3466 = 6'h20 == _myNewVec_11_T_3[5:0] ? myVec_32 : _GEN_3465; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3467 = 6'h21 == _myNewVec_11_T_3[5:0] ? myVec_33 : _GEN_3466; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3468 = 6'h22 == _myNewVec_11_T_3[5:0] ? myVec_34 : _GEN_3467; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3469 = 6'h23 == _myNewVec_11_T_3[5:0] ? myVec_35 : _GEN_3468; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3470 = 6'h24 == _myNewVec_11_T_3[5:0] ? myVec_36 : _GEN_3469; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3471 = 6'h25 == _myNewVec_11_T_3[5:0] ? myVec_37 : _GEN_3470; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3472 = 6'h26 == _myNewVec_11_T_3[5:0] ? myVec_38 : _GEN_3471; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3473 = 6'h27 == _myNewVec_11_T_3[5:0] ? myVec_39 : _GEN_3472; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3474 = 6'h28 == _myNewVec_11_T_3[5:0] ? myVec_40 : _GEN_3473; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3475 = 6'h29 == _myNewVec_11_T_3[5:0] ? myVec_41 : _GEN_3474; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3476 = 6'h2a == _myNewVec_11_T_3[5:0] ? myVec_42 : _GEN_3475; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3477 = 6'h2b == _myNewVec_11_T_3[5:0] ? myVec_43 : _GEN_3476; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3478 = 6'h2c == _myNewVec_11_T_3[5:0] ? myVec_44 : _GEN_3477; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3479 = 6'h2d == _myNewVec_11_T_3[5:0] ? myVec_45 : _GEN_3478; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3480 = 6'h2e == _myNewVec_11_T_3[5:0] ? myVec_46 : _GEN_3479; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3481 = 6'h2f == _myNewVec_11_T_3[5:0] ? myVec_47 : _GEN_3480; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3482 = 6'h30 == _myNewVec_11_T_3[5:0] ? myVec_48 : _GEN_3481; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3483 = 6'h31 == _myNewVec_11_T_3[5:0] ? myVec_49 : _GEN_3482; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3484 = 6'h32 == _myNewVec_11_T_3[5:0] ? myVec_50 : _GEN_3483; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3485 = 6'h33 == _myNewVec_11_T_3[5:0] ? myVec_51 : _GEN_3484; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3486 = 6'h34 == _myNewVec_11_T_3[5:0] ? myVec_52 : _GEN_3485; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3487 = 6'h35 == _myNewVec_11_T_3[5:0] ? myVec_53 : _GEN_3486; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3488 = 6'h36 == _myNewVec_11_T_3[5:0] ? myVec_54 : _GEN_3487; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3489 = 6'h37 == _myNewVec_11_T_3[5:0] ? myVec_55 : _GEN_3488; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3490 = 6'h38 == _myNewVec_11_T_3[5:0] ? myVec_56 : _GEN_3489; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3491 = 6'h39 == _myNewVec_11_T_3[5:0] ? myVec_57 : _GEN_3490; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3492 = 6'h3a == _myNewVec_11_T_3[5:0] ? myVec_58 : _GEN_3491; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3493 = 6'h3b == _myNewVec_11_T_3[5:0] ? myVec_59 : _GEN_3492; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3494 = 6'h3c == _myNewVec_11_T_3[5:0] ? myVec_60 : _GEN_3493; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3495 = 6'h3d == _myNewVec_11_T_3[5:0] ? myVec_61 : _GEN_3494; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3496 = 6'h3e == _myNewVec_11_T_3[5:0] ? myVec_62 : _GEN_3495; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_11 = 6'h3f == _myNewVec_11_T_3[5:0] ? myVec_63 : _GEN_3496; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_10_T_3 = _myNewVec_63_T_1 + 16'h35; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3499 = 6'h1 == _myNewVec_10_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3500 = 6'h2 == _myNewVec_10_T_3[5:0] ? myVec_2 : _GEN_3499; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3501 = 6'h3 == _myNewVec_10_T_3[5:0] ? myVec_3 : _GEN_3500; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3502 = 6'h4 == _myNewVec_10_T_3[5:0] ? myVec_4 : _GEN_3501; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3503 = 6'h5 == _myNewVec_10_T_3[5:0] ? myVec_5 : _GEN_3502; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3504 = 6'h6 == _myNewVec_10_T_3[5:0] ? myVec_6 : _GEN_3503; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3505 = 6'h7 == _myNewVec_10_T_3[5:0] ? myVec_7 : _GEN_3504; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3506 = 6'h8 == _myNewVec_10_T_3[5:0] ? myVec_8 : _GEN_3505; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3507 = 6'h9 == _myNewVec_10_T_3[5:0] ? myVec_9 : _GEN_3506; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3508 = 6'ha == _myNewVec_10_T_3[5:0] ? myVec_10 : _GEN_3507; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3509 = 6'hb == _myNewVec_10_T_3[5:0] ? myVec_11 : _GEN_3508; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3510 = 6'hc == _myNewVec_10_T_3[5:0] ? myVec_12 : _GEN_3509; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3511 = 6'hd == _myNewVec_10_T_3[5:0] ? myVec_13 : _GEN_3510; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3512 = 6'he == _myNewVec_10_T_3[5:0] ? myVec_14 : _GEN_3511; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3513 = 6'hf == _myNewVec_10_T_3[5:0] ? myVec_15 : _GEN_3512; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3514 = 6'h10 == _myNewVec_10_T_3[5:0] ? myVec_16 : _GEN_3513; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3515 = 6'h11 == _myNewVec_10_T_3[5:0] ? myVec_17 : _GEN_3514; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3516 = 6'h12 == _myNewVec_10_T_3[5:0] ? myVec_18 : _GEN_3515; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3517 = 6'h13 == _myNewVec_10_T_3[5:0] ? myVec_19 : _GEN_3516; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3518 = 6'h14 == _myNewVec_10_T_3[5:0] ? myVec_20 : _GEN_3517; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3519 = 6'h15 == _myNewVec_10_T_3[5:0] ? myVec_21 : _GEN_3518; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3520 = 6'h16 == _myNewVec_10_T_3[5:0] ? myVec_22 : _GEN_3519; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3521 = 6'h17 == _myNewVec_10_T_3[5:0] ? myVec_23 : _GEN_3520; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3522 = 6'h18 == _myNewVec_10_T_3[5:0] ? myVec_24 : _GEN_3521; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3523 = 6'h19 == _myNewVec_10_T_3[5:0] ? myVec_25 : _GEN_3522; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3524 = 6'h1a == _myNewVec_10_T_3[5:0] ? myVec_26 : _GEN_3523; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3525 = 6'h1b == _myNewVec_10_T_3[5:0] ? myVec_27 : _GEN_3524; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3526 = 6'h1c == _myNewVec_10_T_3[5:0] ? myVec_28 : _GEN_3525; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3527 = 6'h1d == _myNewVec_10_T_3[5:0] ? myVec_29 : _GEN_3526; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3528 = 6'h1e == _myNewVec_10_T_3[5:0] ? myVec_30 : _GEN_3527; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3529 = 6'h1f == _myNewVec_10_T_3[5:0] ? myVec_31 : _GEN_3528; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3530 = 6'h20 == _myNewVec_10_T_3[5:0] ? myVec_32 : _GEN_3529; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3531 = 6'h21 == _myNewVec_10_T_3[5:0] ? myVec_33 : _GEN_3530; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3532 = 6'h22 == _myNewVec_10_T_3[5:0] ? myVec_34 : _GEN_3531; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3533 = 6'h23 == _myNewVec_10_T_3[5:0] ? myVec_35 : _GEN_3532; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3534 = 6'h24 == _myNewVec_10_T_3[5:0] ? myVec_36 : _GEN_3533; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3535 = 6'h25 == _myNewVec_10_T_3[5:0] ? myVec_37 : _GEN_3534; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3536 = 6'h26 == _myNewVec_10_T_3[5:0] ? myVec_38 : _GEN_3535; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3537 = 6'h27 == _myNewVec_10_T_3[5:0] ? myVec_39 : _GEN_3536; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3538 = 6'h28 == _myNewVec_10_T_3[5:0] ? myVec_40 : _GEN_3537; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3539 = 6'h29 == _myNewVec_10_T_3[5:0] ? myVec_41 : _GEN_3538; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3540 = 6'h2a == _myNewVec_10_T_3[5:0] ? myVec_42 : _GEN_3539; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3541 = 6'h2b == _myNewVec_10_T_3[5:0] ? myVec_43 : _GEN_3540; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3542 = 6'h2c == _myNewVec_10_T_3[5:0] ? myVec_44 : _GEN_3541; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3543 = 6'h2d == _myNewVec_10_T_3[5:0] ? myVec_45 : _GEN_3542; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3544 = 6'h2e == _myNewVec_10_T_3[5:0] ? myVec_46 : _GEN_3543; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3545 = 6'h2f == _myNewVec_10_T_3[5:0] ? myVec_47 : _GEN_3544; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3546 = 6'h30 == _myNewVec_10_T_3[5:0] ? myVec_48 : _GEN_3545; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3547 = 6'h31 == _myNewVec_10_T_3[5:0] ? myVec_49 : _GEN_3546; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3548 = 6'h32 == _myNewVec_10_T_3[5:0] ? myVec_50 : _GEN_3547; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3549 = 6'h33 == _myNewVec_10_T_3[5:0] ? myVec_51 : _GEN_3548; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3550 = 6'h34 == _myNewVec_10_T_3[5:0] ? myVec_52 : _GEN_3549; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3551 = 6'h35 == _myNewVec_10_T_3[5:0] ? myVec_53 : _GEN_3550; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3552 = 6'h36 == _myNewVec_10_T_3[5:0] ? myVec_54 : _GEN_3551; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3553 = 6'h37 == _myNewVec_10_T_3[5:0] ? myVec_55 : _GEN_3552; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3554 = 6'h38 == _myNewVec_10_T_3[5:0] ? myVec_56 : _GEN_3553; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3555 = 6'h39 == _myNewVec_10_T_3[5:0] ? myVec_57 : _GEN_3554; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3556 = 6'h3a == _myNewVec_10_T_3[5:0] ? myVec_58 : _GEN_3555; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3557 = 6'h3b == _myNewVec_10_T_3[5:0] ? myVec_59 : _GEN_3556; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3558 = 6'h3c == _myNewVec_10_T_3[5:0] ? myVec_60 : _GEN_3557; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3559 = 6'h3d == _myNewVec_10_T_3[5:0] ? myVec_61 : _GEN_3558; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3560 = 6'h3e == _myNewVec_10_T_3[5:0] ? myVec_62 : _GEN_3559; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_10 = 6'h3f == _myNewVec_10_T_3[5:0] ? myVec_63 : _GEN_3560; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_9_T_3 = _myNewVec_63_T_1 + 16'h36; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3563 = 6'h1 == _myNewVec_9_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3564 = 6'h2 == _myNewVec_9_T_3[5:0] ? myVec_2 : _GEN_3563; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3565 = 6'h3 == _myNewVec_9_T_3[5:0] ? myVec_3 : _GEN_3564; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3566 = 6'h4 == _myNewVec_9_T_3[5:0] ? myVec_4 : _GEN_3565; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3567 = 6'h5 == _myNewVec_9_T_3[5:0] ? myVec_5 : _GEN_3566; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3568 = 6'h6 == _myNewVec_9_T_3[5:0] ? myVec_6 : _GEN_3567; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3569 = 6'h7 == _myNewVec_9_T_3[5:0] ? myVec_7 : _GEN_3568; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3570 = 6'h8 == _myNewVec_9_T_3[5:0] ? myVec_8 : _GEN_3569; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3571 = 6'h9 == _myNewVec_9_T_3[5:0] ? myVec_9 : _GEN_3570; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3572 = 6'ha == _myNewVec_9_T_3[5:0] ? myVec_10 : _GEN_3571; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3573 = 6'hb == _myNewVec_9_T_3[5:0] ? myVec_11 : _GEN_3572; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3574 = 6'hc == _myNewVec_9_T_3[5:0] ? myVec_12 : _GEN_3573; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3575 = 6'hd == _myNewVec_9_T_3[5:0] ? myVec_13 : _GEN_3574; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3576 = 6'he == _myNewVec_9_T_3[5:0] ? myVec_14 : _GEN_3575; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3577 = 6'hf == _myNewVec_9_T_3[5:0] ? myVec_15 : _GEN_3576; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3578 = 6'h10 == _myNewVec_9_T_3[5:0] ? myVec_16 : _GEN_3577; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3579 = 6'h11 == _myNewVec_9_T_3[5:0] ? myVec_17 : _GEN_3578; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3580 = 6'h12 == _myNewVec_9_T_3[5:0] ? myVec_18 : _GEN_3579; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3581 = 6'h13 == _myNewVec_9_T_3[5:0] ? myVec_19 : _GEN_3580; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3582 = 6'h14 == _myNewVec_9_T_3[5:0] ? myVec_20 : _GEN_3581; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3583 = 6'h15 == _myNewVec_9_T_3[5:0] ? myVec_21 : _GEN_3582; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3584 = 6'h16 == _myNewVec_9_T_3[5:0] ? myVec_22 : _GEN_3583; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3585 = 6'h17 == _myNewVec_9_T_3[5:0] ? myVec_23 : _GEN_3584; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3586 = 6'h18 == _myNewVec_9_T_3[5:0] ? myVec_24 : _GEN_3585; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3587 = 6'h19 == _myNewVec_9_T_3[5:0] ? myVec_25 : _GEN_3586; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3588 = 6'h1a == _myNewVec_9_T_3[5:0] ? myVec_26 : _GEN_3587; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3589 = 6'h1b == _myNewVec_9_T_3[5:0] ? myVec_27 : _GEN_3588; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3590 = 6'h1c == _myNewVec_9_T_3[5:0] ? myVec_28 : _GEN_3589; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3591 = 6'h1d == _myNewVec_9_T_3[5:0] ? myVec_29 : _GEN_3590; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3592 = 6'h1e == _myNewVec_9_T_3[5:0] ? myVec_30 : _GEN_3591; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3593 = 6'h1f == _myNewVec_9_T_3[5:0] ? myVec_31 : _GEN_3592; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3594 = 6'h20 == _myNewVec_9_T_3[5:0] ? myVec_32 : _GEN_3593; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3595 = 6'h21 == _myNewVec_9_T_3[5:0] ? myVec_33 : _GEN_3594; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3596 = 6'h22 == _myNewVec_9_T_3[5:0] ? myVec_34 : _GEN_3595; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3597 = 6'h23 == _myNewVec_9_T_3[5:0] ? myVec_35 : _GEN_3596; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3598 = 6'h24 == _myNewVec_9_T_3[5:0] ? myVec_36 : _GEN_3597; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3599 = 6'h25 == _myNewVec_9_T_3[5:0] ? myVec_37 : _GEN_3598; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3600 = 6'h26 == _myNewVec_9_T_3[5:0] ? myVec_38 : _GEN_3599; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3601 = 6'h27 == _myNewVec_9_T_3[5:0] ? myVec_39 : _GEN_3600; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3602 = 6'h28 == _myNewVec_9_T_3[5:0] ? myVec_40 : _GEN_3601; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3603 = 6'h29 == _myNewVec_9_T_3[5:0] ? myVec_41 : _GEN_3602; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3604 = 6'h2a == _myNewVec_9_T_3[5:0] ? myVec_42 : _GEN_3603; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3605 = 6'h2b == _myNewVec_9_T_3[5:0] ? myVec_43 : _GEN_3604; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3606 = 6'h2c == _myNewVec_9_T_3[5:0] ? myVec_44 : _GEN_3605; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3607 = 6'h2d == _myNewVec_9_T_3[5:0] ? myVec_45 : _GEN_3606; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3608 = 6'h2e == _myNewVec_9_T_3[5:0] ? myVec_46 : _GEN_3607; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3609 = 6'h2f == _myNewVec_9_T_3[5:0] ? myVec_47 : _GEN_3608; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3610 = 6'h30 == _myNewVec_9_T_3[5:0] ? myVec_48 : _GEN_3609; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3611 = 6'h31 == _myNewVec_9_T_3[5:0] ? myVec_49 : _GEN_3610; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3612 = 6'h32 == _myNewVec_9_T_3[5:0] ? myVec_50 : _GEN_3611; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3613 = 6'h33 == _myNewVec_9_T_3[5:0] ? myVec_51 : _GEN_3612; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3614 = 6'h34 == _myNewVec_9_T_3[5:0] ? myVec_52 : _GEN_3613; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3615 = 6'h35 == _myNewVec_9_T_3[5:0] ? myVec_53 : _GEN_3614; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3616 = 6'h36 == _myNewVec_9_T_3[5:0] ? myVec_54 : _GEN_3615; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3617 = 6'h37 == _myNewVec_9_T_3[5:0] ? myVec_55 : _GEN_3616; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3618 = 6'h38 == _myNewVec_9_T_3[5:0] ? myVec_56 : _GEN_3617; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3619 = 6'h39 == _myNewVec_9_T_3[5:0] ? myVec_57 : _GEN_3618; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3620 = 6'h3a == _myNewVec_9_T_3[5:0] ? myVec_58 : _GEN_3619; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3621 = 6'h3b == _myNewVec_9_T_3[5:0] ? myVec_59 : _GEN_3620; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3622 = 6'h3c == _myNewVec_9_T_3[5:0] ? myVec_60 : _GEN_3621; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3623 = 6'h3d == _myNewVec_9_T_3[5:0] ? myVec_61 : _GEN_3622; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3624 = 6'h3e == _myNewVec_9_T_3[5:0] ? myVec_62 : _GEN_3623; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_9 = 6'h3f == _myNewVec_9_T_3[5:0] ? myVec_63 : _GEN_3624; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_8_T_3 = _myNewVec_63_T_1 + 16'h37; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3627 = 6'h1 == _myNewVec_8_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3628 = 6'h2 == _myNewVec_8_T_3[5:0] ? myVec_2 : _GEN_3627; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3629 = 6'h3 == _myNewVec_8_T_3[5:0] ? myVec_3 : _GEN_3628; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3630 = 6'h4 == _myNewVec_8_T_3[5:0] ? myVec_4 : _GEN_3629; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3631 = 6'h5 == _myNewVec_8_T_3[5:0] ? myVec_5 : _GEN_3630; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3632 = 6'h6 == _myNewVec_8_T_3[5:0] ? myVec_6 : _GEN_3631; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3633 = 6'h7 == _myNewVec_8_T_3[5:0] ? myVec_7 : _GEN_3632; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3634 = 6'h8 == _myNewVec_8_T_3[5:0] ? myVec_8 : _GEN_3633; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3635 = 6'h9 == _myNewVec_8_T_3[5:0] ? myVec_9 : _GEN_3634; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3636 = 6'ha == _myNewVec_8_T_3[5:0] ? myVec_10 : _GEN_3635; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3637 = 6'hb == _myNewVec_8_T_3[5:0] ? myVec_11 : _GEN_3636; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3638 = 6'hc == _myNewVec_8_T_3[5:0] ? myVec_12 : _GEN_3637; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3639 = 6'hd == _myNewVec_8_T_3[5:0] ? myVec_13 : _GEN_3638; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3640 = 6'he == _myNewVec_8_T_3[5:0] ? myVec_14 : _GEN_3639; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3641 = 6'hf == _myNewVec_8_T_3[5:0] ? myVec_15 : _GEN_3640; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3642 = 6'h10 == _myNewVec_8_T_3[5:0] ? myVec_16 : _GEN_3641; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3643 = 6'h11 == _myNewVec_8_T_3[5:0] ? myVec_17 : _GEN_3642; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3644 = 6'h12 == _myNewVec_8_T_3[5:0] ? myVec_18 : _GEN_3643; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3645 = 6'h13 == _myNewVec_8_T_3[5:0] ? myVec_19 : _GEN_3644; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3646 = 6'h14 == _myNewVec_8_T_3[5:0] ? myVec_20 : _GEN_3645; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3647 = 6'h15 == _myNewVec_8_T_3[5:0] ? myVec_21 : _GEN_3646; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3648 = 6'h16 == _myNewVec_8_T_3[5:0] ? myVec_22 : _GEN_3647; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3649 = 6'h17 == _myNewVec_8_T_3[5:0] ? myVec_23 : _GEN_3648; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3650 = 6'h18 == _myNewVec_8_T_3[5:0] ? myVec_24 : _GEN_3649; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3651 = 6'h19 == _myNewVec_8_T_3[5:0] ? myVec_25 : _GEN_3650; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3652 = 6'h1a == _myNewVec_8_T_3[5:0] ? myVec_26 : _GEN_3651; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3653 = 6'h1b == _myNewVec_8_T_3[5:0] ? myVec_27 : _GEN_3652; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3654 = 6'h1c == _myNewVec_8_T_3[5:0] ? myVec_28 : _GEN_3653; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3655 = 6'h1d == _myNewVec_8_T_3[5:0] ? myVec_29 : _GEN_3654; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3656 = 6'h1e == _myNewVec_8_T_3[5:0] ? myVec_30 : _GEN_3655; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3657 = 6'h1f == _myNewVec_8_T_3[5:0] ? myVec_31 : _GEN_3656; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3658 = 6'h20 == _myNewVec_8_T_3[5:0] ? myVec_32 : _GEN_3657; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3659 = 6'h21 == _myNewVec_8_T_3[5:0] ? myVec_33 : _GEN_3658; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3660 = 6'h22 == _myNewVec_8_T_3[5:0] ? myVec_34 : _GEN_3659; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3661 = 6'h23 == _myNewVec_8_T_3[5:0] ? myVec_35 : _GEN_3660; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3662 = 6'h24 == _myNewVec_8_T_3[5:0] ? myVec_36 : _GEN_3661; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3663 = 6'h25 == _myNewVec_8_T_3[5:0] ? myVec_37 : _GEN_3662; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3664 = 6'h26 == _myNewVec_8_T_3[5:0] ? myVec_38 : _GEN_3663; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3665 = 6'h27 == _myNewVec_8_T_3[5:0] ? myVec_39 : _GEN_3664; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3666 = 6'h28 == _myNewVec_8_T_3[5:0] ? myVec_40 : _GEN_3665; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3667 = 6'h29 == _myNewVec_8_T_3[5:0] ? myVec_41 : _GEN_3666; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3668 = 6'h2a == _myNewVec_8_T_3[5:0] ? myVec_42 : _GEN_3667; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3669 = 6'h2b == _myNewVec_8_T_3[5:0] ? myVec_43 : _GEN_3668; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3670 = 6'h2c == _myNewVec_8_T_3[5:0] ? myVec_44 : _GEN_3669; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3671 = 6'h2d == _myNewVec_8_T_3[5:0] ? myVec_45 : _GEN_3670; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3672 = 6'h2e == _myNewVec_8_T_3[5:0] ? myVec_46 : _GEN_3671; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3673 = 6'h2f == _myNewVec_8_T_3[5:0] ? myVec_47 : _GEN_3672; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3674 = 6'h30 == _myNewVec_8_T_3[5:0] ? myVec_48 : _GEN_3673; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3675 = 6'h31 == _myNewVec_8_T_3[5:0] ? myVec_49 : _GEN_3674; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3676 = 6'h32 == _myNewVec_8_T_3[5:0] ? myVec_50 : _GEN_3675; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3677 = 6'h33 == _myNewVec_8_T_3[5:0] ? myVec_51 : _GEN_3676; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3678 = 6'h34 == _myNewVec_8_T_3[5:0] ? myVec_52 : _GEN_3677; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3679 = 6'h35 == _myNewVec_8_T_3[5:0] ? myVec_53 : _GEN_3678; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3680 = 6'h36 == _myNewVec_8_T_3[5:0] ? myVec_54 : _GEN_3679; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3681 = 6'h37 == _myNewVec_8_T_3[5:0] ? myVec_55 : _GEN_3680; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3682 = 6'h38 == _myNewVec_8_T_3[5:0] ? myVec_56 : _GEN_3681; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3683 = 6'h39 == _myNewVec_8_T_3[5:0] ? myVec_57 : _GEN_3682; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3684 = 6'h3a == _myNewVec_8_T_3[5:0] ? myVec_58 : _GEN_3683; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3685 = 6'h3b == _myNewVec_8_T_3[5:0] ? myVec_59 : _GEN_3684; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3686 = 6'h3c == _myNewVec_8_T_3[5:0] ? myVec_60 : _GEN_3685; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3687 = 6'h3d == _myNewVec_8_T_3[5:0] ? myVec_61 : _GEN_3686; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3688 = 6'h3e == _myNewVec_8_T_3[5:0] ? myVec_62 : _GEN_3687; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_8 = 6'h3f == _myNewVec_8_T_3[5:0] ? myVec_63 : _GEN_3688; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_7_T_3 = _myNewVec_63_T_1 + 16'h38; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3691 = 6'h1 == _myNewVec_7_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3692 = 6'h2 == _myNewVec_7_T_3[5:0] ? myVec_2 : _GEN_3691; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3693 = 6'h3 == _myNewVec_7_T_3[5:0] ? myVec_3 : _GEN_3692; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3694 = 6'h4 == _myNewVec_7_T_3[5:0] ? myVec_4 : _GEN_3693; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3695 = 6'h5 == _myNewVec_7_T_3[5:0] ? myVec_5 : _GEN_3694; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3696 = 6'h6 == _myNewVec_7_T_3[5:0] ? myVec_6 : _GEN_3695; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3697 = 6'h7 == _myNewVec_7_T_3[5:0] ? myVec_7 : _GEN_3696; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3698 = 6'h8 == _myNewVec_7_T_3[5:0] ? myVec_8 : _GEN_3697; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3699 = 6'h9 == _myNewVec_7_T_3[5:0] ? myVec_9 : _GEN_3698; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3700 = 6'ha == _myNewVec_7_T_3[5:0] ? myVec_10 : _GEN_3699; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3701 = 6'hb == _myNewVec_7_T_3[5:0] ? myVec_11 : _GEN_3700; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3702 = 6'hc == _myNewVec_7_T_3[5:0] ? myVec_12 : _GEN_3701; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3703 = 6'hd == _myNewVec_7_T_3[5:0] ? myVec_13 : _GEN_3702; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3704 = 6'he == _myNewVec_7_T_3[5:0] ? myVec_14 : _GEN_3703; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3705 = 6'hf == _myNewVec_7_T_3[5:0] ? myVec_15 : _GEN_3704; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3706 = 6'h10 == _myNewVec_7_T_3[5:0] ? myVec_16 : _GEN_3705; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3707 = 6'h11 == _myNewVec_7_T_3[5:0] ? myVec_17 : _GEN_3706; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3708 = 6'h12 == _myNewVec_7_T_3[5:0] ? myVec_18 : _GEN_3707; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3709 = 6'h13 == _myNewVec_7_T_3[5:0] ? myVec_19 : _GEN_3708; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3710 = 6'h14 == _myNewVec_7_T_3[5:0] ? myVec_20 : _GEN_3709; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3711 = 6'h15 == _myNewVec_7_T_3[5:0] ? myVec_21 : _GEN_3710; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3712 = 6'h16 == _myNewVec_7_T_3[5:0] ? myVec_22 : _GEN_3711; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3713 = 6'h17 == _myNewVec_7_T_3[5:0] ? myVec_23 : _GEN_3712; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3714 = 6'h18 == _myNewVec_7_T_3[5:0] ? myVec_24 : _GEN_3713; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3715 = 6'h19 == _myNewVec_7_T_3[5:0] ? myVec_25 : _GEN_3714; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3716 = 6'h1a == _myNewVec_7_T_3[5:0] ? myVec_26 : _GEN_3715; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3717 = 6'h1b == _myNewVec_7_T_3[5:0] ? myVec_27 : _GEN_3716; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3718 = 6'h1c == _myNewVec_7_T_3[5:0] ? myVec_28 : _GEN_3717; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3719 = 6'h1d == _myNewVec_7_T_3[5:0] ? myVec_29 : _GEN_3718; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3720 = 6'h1e == _myNewVec_7_T_3[5:0] ? myVec_30 : _GEN_3719; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3721 = 6'h1f == _myNewVec_7_T_3[5:0] ? myVec_31 : _GEN_3720; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3722 = 6'h20 == _myNewVec_7_T_3[5:0] ? myVec_32 : _GEN_3721; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3723 = 6'h21 == _myNewVec_7_T_3[5:0] ? myVec_33 : _GEN_3722; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3724 = 6'h22 == _myNewVec_7_T_3[5:0] ? myVec_34 : _GEN_3723; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3725 = 6'h23 == _myNewVec_7_T_3[5:0] ? myVec_35 : _GEN_3724; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3726 = 6'h24 == _myNewVec_7_T_3[5:0] ? myVec_36 : _GEN_3725; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3727 = 6'h25 == _myNewVec_7_T_3[5:0] ? myVec_37 : _GEN_3726; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3728 = 6'h26 == _myNewVec_7_T_3[5:0] ? myVec_38 : _GEN_3727; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3729 = 6'h27 == _myNewVec_7_T_3[5:0] ? myVec_39 : _GEN_3728; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3730 = 6'h28 == _myNewVec_7_T_3[5:0] ? myVec_40 : _GEN_3729; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3731 = 6'h29 == _myNewVec_7_T_3[5:0] ? myVec_41 : _GEN_3730; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3732 = 6'h2a == _myNewVec_7_T_3[5:0] ? myVec_42 : _GEN_3731; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3733 = 6'h2b == _myNewVec_7_T_3[5:0] ? myVec_43 : _GEN_3732; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3734 = 6'h2c == _myNewVec_7_T_3[5:0] ? myVec_44 : _GEN_3733; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3735 = 6'h2d == _myNewVec_7_T_3[5:0] ? myVec_45 : _GEN_3734; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3736 = 6'h2e == _myNewVec_7_T_3[5:0] ? myVec_46 : _GEN_3735; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3737 = 6'h2f == _myNewVec_7_T_3[5:0] ? myVec_47 : _GEN_3736; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3738 = 6'h30 == _myNewVec_7_T_3[5:0] ? myVec_48 : _GEN_3737; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3739 = 6'h31 == _myNewVec_7_T_3[5:0] ? myVec_49 : _GEN_3738; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3740 = 6'h32 == _myNewVec_7_T_3[5:0] ? myVec_50 : _GEN_3739; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3741 = 6'h33 == _myNewVec_7_T_3[5:0] ? myVec_51 : _GEN_3740; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3742 = 6'h34 == _myNewVec_7_T_3[5:0] ? myVec_52 : _GEN_3741; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3743 = 6'h35 == _myNewVec_7_T_3[5:0] ? myVec_53 : _GEN_3742; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3744 = 6'h36 == _myNewVec_7_T_3[5:0] ? myVec_54 : _GEN_3743; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3745 = 6'h37 == _myNewVec_7_T_3[5:0] ? myVec_55 : _GEN_3744; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3746 = 6'h38 == _myNewVec_7_T_3[5:0] ? myVec_56 : _GEN_3745; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3747 = 6'h39 == _myNewVec_7_T_3[5:0] ? myVec_57 : _GEN_3746; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3748 = 6'h3a == _myNewVec_7_T_3[5:0] ? myVec_58 : _GEN_3747; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3749 = 6'h3b == _myNewVec_7_T_3[5:0] ? myVec_59 : _GEN_3748; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3750 = 6'h3c == _myNewVec_7_T_3[5:0] ? myVec_60 : _GEN_3749; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3751 = 6'h3d == _myNewVec_7_T_3[5:0] ? myVec_61 : _GEN_3750; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3752 = 6'h3e == _myNewVec_7_T_3[5:0] ? myVec_62 : _GEN_3751; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_7 = 6'h3f == _myNewVec_7_T_3[5:0] ? myVec_63 : _GEN_3752; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_6_T_3 = _myNewVec_63_T_1 + 16'h39; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3755 = 6'h1 == _myNewVec_6_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3756 = 6'h2 == _myNewVec_6_T_3[5:0] ? myVec_2 : _GEN_3755; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3757 = 6'h3 == _myNewVec_6_T_3[5:0] ? myVec_3 : _GEN_3756; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3758 = 6'h4 == _myNewVec_6_T_3[5:0] ? myVec_4 : _GEN_3757; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3759 = 6'h5 == _myNewVec_6_T_3[5:0] ? myVec_5 : _GEN_3758; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3760 = 6'h6 == _myNewVec_6_T_3[5:0] ? myVec_6 : _GEN_3759; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3761 = 6'h7 == _myNewVec_6_T_3[5:0] ? myVec_7 : _GEN_3760; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3762 = 6'h8 == _myNewVec_6_T_3[5:0] ? myVec_8 : _GEN_3761; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3763 = 6'h9 == _myNewVec_6_T_3[5:0] ? myVec_9 : _GEN_3762; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3764 = 6'ha == _myNewVec_6_T_3[5:0] ? myVec_10 : _GEN_3763; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3765 = 6'hb == _myNewVec_6_T_3[5:0] ? myVec_11 : _GEN_3764; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3766 = 6'hc == _myNewVec_6_T_3[5:0] ? myVec_12 : _GEN_3765; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3767 = 6'hd == _myNewVec_6_T_3[5:0] ? myVec_13 : _GEN_3766; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3768 = 6'he == _myNewVec_6_T_3[5:0] ? myVec_14 : _GEN_3767; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3769 = 6'hf == _myNewVec_6_T_3[5:0] ? myVec_15 : _GEN_3768; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3770 = 6'h10 == _myNewVec_6_T_3[5:0] ? myVec_16 : _GEN_3769; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3771 = 6'h11 == _myNewVec_6_T_3[5:0] ? myVec_17 : _GEN_3770; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3772 = 6'h12 == _myNewVec_6_T_3[5:0] ? myVec_18 : _GEN_3771; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3773 = 6'h13 == _myNewVec_6_T_3[5:0] ? myVec_19 : _GEN_3772; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3774 = 6'h14 == _myNewVec_6_T_3[5:0] ? myVec_20 : _GEN_3773; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3775 = 6'h15 == _myNewVec_6_T_3[5:0] ? myVec_21 : _GEN_3774; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3776 = 6'h16 == _myNewVec_6_T_3[5:0] ? myVec_22 : _GEN_3775; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3777 = 6'h17 == _myNewVec_6_T_3[5:0] ? myVec_23 : _GEN_3776; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3778 = 6'h18 == _myNewVec_6_T_3[5:0] ? myVec_24 : _GEN_3777; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3779 = 6'h19 == _myNewVec_6_T_3[5:0] ? myVec_25 : _GEN_3778; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3780 = 6'h1a == _myNewVec_6_T_3[5:0] ? myVec_26 : _GEN_3779; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3781 = 6'h1b == _myNewVec_6_T_3[5:0] ? myVec_27 : _GEN_3780; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3782 = 6'h1c == _myNewVec_6_T_3[5:0] ? myVec_28 : _GEN_3781; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3783 = 6'h1d == _myNewVec_6_T_3[5:0] ? myVec_29 : _GEN_3782; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3784 = 6'h1e == _myNewVec_6_T_3[5:0] ? myVec_30 : _GEN_3783; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3785 = 6'h1f == _myNewVec_6_T_3[5:0] ? myVec_31 : _GEN_3784; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3786 = 6'h20 == _myNewVec_6_T_3[5:0] ? myVec_32 : _GEN_3785; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3787 = 6'h21 == _myNewVec_6_T_3[5:0] ? myVec_33 : _GEN_3786; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3788 = 6'h22 == _myNewVec_6_T_3[5:0] ? myVec_34 : _GEN_3787; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3789 = 6'h23 == _myNewVec_6_T_3[5:0] ? myVec_35 : _GEN_3788; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3790 = 6'h24 == _myNewVec_6_T_3[5:0] ? myVec_36 : _GEN_3789; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3791 = 6'h25 == _myNewVec_6_T_3[5:0] ? myVec_37 : _GEN_3790; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3792 = 6'h26 == _myNewVec_6_T_3[5:0] ? myVec_38 : _GEN_3791; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3793 = 6'h27 == _myNewVec_6_T_3[5:0] ? myVec_39 : _GEN_3792; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3794 = 6'h28 == _myNewVec_6_T_3[5:0] ? myVec_40 : _GEN_3793; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3795 = 6'h29 == _myNewVec_6_T_3[5:0] ? myVec_41 : _GEN_3794; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3796 = 6'h2a == _myNewVec_6_T_3[5:0] ? myVec_42 : _GEN_3795; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3797 = 6'h2b == _myNewVec_6_T_3[5:0] ? myVec_43 : _GEN_3796; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3798 = 6'h2c == _myNewVec_6_T_3[5:0] ? myVec_44 : _GEN_3797; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3799 = 6'h2d == _myNewVec_6_T_3[5:0] ? myVec_45 : _GEN_3798; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3800 = 6'h2e == _myNewVec_6_T_3[5:0] ? myVec_46 : _GEN_3799; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3801 = 6'h2f == _myNewVec_6_T_3[5:0] ? myVec_47 : _GEN_3800; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3802 = 6'h30 == _myNewVec_6_T_3[5:0] ? myVec_48 : _GEN_3801; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3803 = 6'h31 == _myNewVec_6_T_3[5:0] ? myVec_49 : _GEN_3802; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3804 = 6'h32 == _myNewVec_6_T_3[5:0] ? myVec_50 : _GEN_3803; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3805 = 6'h33 == _myNewVec_6_T_3[5:0] ? myVec_51 : _GEN_3804; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3806 = 6'h34 == _myNewVec_6_T_3[5:0] ? myVec_52 : _GEN_3805; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3807 = 6'h35 == _myNewVec_6_T_3[5:0] ? myVec_53 : _GEN_3806; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3808 = 6'h36 == _myNewVec_6_T_3[5:0] ? myVec_54 : _GEN_3807; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3809 = 6'h37 == _myNewVec_6_T_3[5:0] ? myVec_55 : _GEN_3808; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3810 = 6'h38 == _myNewVec_6_T_3[5:0] ? myVec_56 : _GEN_3809; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3811 = 6'h39 == _myNewVec_6_T_3[5:0] ? myVec_57 : _GEN_3810; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3812 = 6'h3a == _myNewVec_6_T_3[5:0] ? myVec_58 : _GEN_3811; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3813 = 6'h3b == _myNewVec_6_T_3[5:0] ? myVec_59 : _GEN_3812; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3814 = 6'h3c == _myNewVec_6_T_3[5:0] ? myVec_60 : _GEN_3813; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3815 = 6'h3d == _myNewVec_6_T_3[5:0] ? myVec_61 : _GEN_3814; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3816 = 6'h3e == _myNewVec_6_T_3[5:0] ? myVec_62 : _GEN_3815; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_6 = 6'h3f == _myNewVec_6_T_3[5:0] ? myVec_63 : _GEN_3816; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_5_T_3 = _myNewVec_63_T_1 + 16'h3a; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3819 = 6'h1 == _myNewVec_5_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3820 = 6'h2 == _myNewVec_5_T_3[5:0] ? myVec_2 : _GEN_3819; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3821 = 6'h3 == _myNewVec_5_T_3[5:0] ? myVec_3 : _GEN_3820; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3822 = 6'h4 == _myNewVec_5_T_3[5:0] ? myVec_4 : _GEN_3821; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3823 = 6'h5 == _myNewVec_5_T_3[5:0] ? myVec_5 : _GEN_3822; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3824 = 6'h6 == _myNewVec_5_T_3[5:0] ? myVec_6 : _GEN_3823; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3825 = 6'h7 == _myNewVec_5_T_3[5:0] ? myVec_7 : _GEN_3824; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3826 = 6'h8 == _myNewVec_5_T_3[5:0] ? myVec_8 : _GEN_3825; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3827 = 6'h9 == _myNewVec_5_T_3[5:0] ? myVec_9 : _GEN_3826; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3828 = 6'ha == _myNewVec_5_T_3[5:0] ? myVec_10 : _GEN_3827; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3829 = 6'hb == _myNewVec_5_T_3[5:0] ? myVec_11 : _GEN_3828; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3830 = 6'hc == _myNewVec_5_T_3[5:0] ? myVec_12 : _GEN_3829; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3831 = 6'hd == _myNewVec_5_T_3[5:0] ? myVec_13 : _GEN_3830; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3832 = 6'he == _myNewVec_5_T_3[5:0] ? myVec_14 : _GEN_3831; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3833 = 6'hf == _myNewVec_5_T_3[5:0] ? myVec_15 : _GEN_3832; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3834 = 6'h10 == _myNewVec_5_T_3[5:0] ? myVec_16 : _GEN_3833; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3835 = 6'h11 == _myNewVec_5_T_3[5:0] ? myVec_17 : _GEN_3834; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3836 = 6'h12 == _myNewVec_5_T_3[5:0] ? myVec_18 : _GEN_3835; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3837 = 6'h13 == _myNewVec_5_T_3[5:0] ? myVec_19 : _GEN_3836; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3838 = 6'h14 == _myNewVec_5_T_3[5:0] ? myVec_20 : _GEN_3837; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3839 = 6'h15 == _myNewVec_5_T_3[5:0] ? myVec_21 : _GEN_3838; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3840 = 6'h16 == _myNewVec_5_T_3[5:0] ? myVec_22 : _GEN_3839; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3841 = 6'h17 == _myNewVec_5_T_3[5:0] ? myVec_23 : _GEN_3840; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3842 = 6'h18 == _myNewVec_5_T_3[5:0] ? myVec_24 : _GEN_3841; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3843 = 6'h19 == _myNewVec_5_T_3[5:0] ? myVec_25 : _GEN_3842; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3844 = 6'h1a == _myNewVec_5_T_3[5:0] ? myVec_26 : _GEN_3843; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3845 = 6'h1b == _myNewVec_5_T_3[5:0] ? myVec_27 : _GEN_3844; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3846 = 6'h1c == _myNewVec_5_T_3[5:0] ? myVec_28 : _GEN_3845; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3847 = 6'h1d == _myNewVec_5_T_3[5:0] ? myVec_29 : _GEN_3846; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3848 = 6'h1e == _myNewVec_5_T_3[5:0] ? myVec_30 : _GEN_3847; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3849 = 6'h1f == _myNewVec_5_T_3[5:0] ? myVec_31 : _GEN_3848; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3850 = 6'h20 == _myNewVec_5_T_3[5:0] ? myVec_32 : _GEN_3849; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3851 = 6'h21 == _myNewVec_5_T_3[5:0] ? myVec_33 : _GEN_3850; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3852 = 6'h22 == _myNewVec_5_T_3[5:0] ? myVec_34 : _GEN_3851; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3853 = 6'h23 == _myNewVec_5_T_3[5:0] ? myVec_35 : _GEN_3852; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3854 = 6'h24 == _myNewVec_5_T_3[5:0] ? myVec_36 : _GEN_3853; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3855 = 6'h25 == _myNewVec_5_T_3[5:0] ? myVec_37 : _GEN_3854; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3856 = 6'h26 == _myNewVec_5_T_3[5:0] ? myVec_38 : _GEN_3855; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3857 = 6'h27 == _myNewVec_5_T_3[5:0] ? myVec_39 : _GEN_3856; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3858 = 6'h28 == _myNewVec_5_T_3[5:0] ? myVec_40 : _GEN_3857; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3859 = 6'h29 == _myNewVec_5_T_3[5:0] ? myVec_41 : _GEN_3858; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3860 = 6'h2a == _myNewVec_5_T_3[5:0] ? myVec_42 : _GEN_3859; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3861 = 6'h2b == _myNewVec_5_T_3[5:0] ? myVec_43 : _GEN_3860; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3862 = 6'h2c == _myNewVec_5_T_3[5:0] ? myVec_44 : _GEN_3861; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3863 = 6'h2d == _myNewVec_5_T_3[5:0] ? myVec_45 : _GEN_3862; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3864 = 6'h2e == _myNewVec_5_T_3[5:0] ? myVec_46 : _GEN_3863; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3865 = 6'h2f == _myNewVec_5_T_3[5:0] ? myVec_47 : _GEN_3864; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3866 = 6'h30 == _myNewVec_5_T_3[5:0] ? myVec_48 : _GEN_3865; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3867 = 6'h31 == _myNewVec_5_T_3[5:0] ? myVec_49 : _GEN_3866; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3868 = 6'h32 == _myNewVec_5_T_3[5:0] ? myVec_50 : _GEN_3867; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3869 = 6'h33 == _myNewVec_5_T_3[5:0] ? myVec_51 : _GEN_3868; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3870 = 6'h34 == _myNewVec_5_T_3[5:0] ? myVec_52 : _GEN_3869; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3871 = 6'h35 == _myNewVec_5_T_3[5:0] ? myVec_53 : _GEN_3870; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3872 = 6'h36 == _myNewVec_5_T_3[5:0] ? myVec_54 : _GEN_3871; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3873 = 6'h37 == _myNewVec_5_T_3[5:0] ? myVec_55 : _GEN_3872; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3874 = 6'h38 == _myNewVec_5_T_3[5:0] ? myVec_56 : _GEN_3873; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3875 = 6'h39 == _myNewVec_5_T_3[5:0] ? myVec_57 : _GEN_3874; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3876 = 6'h3a == _myNewVec_5_T_3[5:0] ? myVec_58 : _GEN_3875; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3877 = 6'h3b == _myNewVec_5_T_3[5:0] ? myVec_59 : _GEN_3876; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3878 = 6'h3c == _myNewVec_5_T_3[5:0] ? myVec_60 : _GEN_3877; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3879 = 6'h3d == _myNewVec_5_T_3[5:0] ? myVec_61 : _GEN_3878; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3880 = 6'h3e == _myNewVec_5_T_3[5:0] ? myVec_62 : _GEN_3879; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_5 = 6'h3f == _myNewVec_5_T_3[5:0] ? myVec_63 : _GEN_3880; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_4_T_3 = _myNewVec_63_T_1 + 16'h3b; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3883 = 6'h1 == _myNewVec_4_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3884 = 6'h2 == _myNewVec_4_T_3[5:0] ? myVec_2 : _GEN_3883; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3885 = 6'h3 == _myNewVec_4_T_3[5:0] ? myVec_3 : _GEN_3884; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3886 = 6'h4 == _myNewVec_4_T_3[5:0] ? myVec_4 : _GEN_3885; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3887 = 6'h5 == _myNewVec_4_T_3[5:0] ? myVec_5 : _GEN_3886; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3888 = 6'h6 == _myNewVec_4_T_3[5:0] ? myVec_6 : _GEN_3887; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3889 = 6'h7 == _myNewVec_4_T_3[5:0] ? myVec_7 : _GEN_3888; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3890 = 6'h8 == _myNewVec_4_T_3[5:0] ? myVec_8 : _GEN_3889; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3891 = 6'h9 == _myNewVec_4_T_3[5:0] ? myVec_9 : _GEN_3890; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3892 = 6'ha == _myNewVec_4_T_3[5:0] ? myVec_10 : _GEN_3891; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3893 = 6'hb == _myNewVec_4_T_3[5:0] ? myVec_11 : _GEN_3892; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3894 = 6'hc == _myNewVec_4_T_3[5:0] ? myVec_12 : _GEN_3893; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3895 = 6'hd == _myNewVec_4_T_3[5:0] ? myVec_13 : _GEN_3894; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3896 = 6'he == _myNewVec_4_T_3[5:0] ? myVec_14 : _GEN_3895; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3897 = 6'hf == _myNewVec_4_T_3[5:0] ? myVec_15 : _GEN_3896; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3898 = 6'h10 == _myNewVec_4_T_3[5:0] ? myVec_16 : _GEN_3897; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3899 = 6'h11 == _myNewVec_4_T_3[5:0] ? myVec_17 : _GEN_3898; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3900 = 6'h12 == _myNewVec_4_T_3[5:0] ? myVec_18 : _GEN_3899; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3901 = 6'h13 == _myNewVec_4_T_3[5:0] ? myVec_19 : _GEN_3900; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3902 = 6'h14 == _myNewVec_4_T_3[5:0] ? myVec_20 : _GEN_3901; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3903 = 6'h15 == _myNewVec_4_T_3[5:0] ? myVec_21 : _GEN_3902; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3904 = 6'h16 == _myNewVec_4_T_3[5:0] ? myVec_22 : _GEN_3903; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3905 = 6'h17 == _myNewVec_4_T_3[5:0] ? myVec_23 : _GEN_3904; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3906 = 6'h18 == _myNewVec_4_T_3[5:0] ? myVec_24 : _GEN_3905; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3907 = 6'h19 == _myNewVec_4_T_3[5:0] ? myVec_25 : _GEN_3906; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3908 = 6'h1a == _myNewVec_4_T_3[5:0] ? myVec_26 : _GEN_3907; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3909 = 6'h1b == _myNewVec_4_T_3[5:0] ? myVec_27 : _GEN_3908; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3910 = 6'h1c == _myNewVec_4_T_3[5:0] ? myVec_28 : _GEN_3909; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3911 = 6'h1d == _myNewVec_4_T_3[5:0] ? myVec_29 : _GEN_3910; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3912 = 6'h1e == _myNewVec_4_T_3[5:0] ? myVec_30 : _GEN_3911; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3913 = 6'h1f == _myNewVec_4_T_3[5:0] ? myVec_31 : _GEN_3912; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3914 = 6'h20 == _myNewVec_4_T_3[5:0] ? myVec_32 : _GEN_3913; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3915 = 6'h21 == _myNewVec_4_T_3[5:0] ? myVec_33 : _GEN_3914; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3916 = 6'h22 == _myNewVec_4_T_3[5:0] ? myVec_34 : _GEN_3915; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3917 = 6'h23 == _myNewVec_4_T_3[5:0] ? myVec_35 : _GEN_3916; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3918 = 6'h24 == _myNewVec_4_T_3[5:0] ? myVec_36 : _GEN_3917; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3919 = 6'h25 == _myNewVec_4_T_3[5:0] ? myVec_37 : _GEN_3918; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3920 = 6'h26 == _myNewVec_4_T_3[5:0] ? myVec_38 : _GEN_3919; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3921 = 6'h27 == _myNewVec_4_T_3[5:0] ? myVec_39 : _GEN_3920; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3922 = 6'h28 == _myNewVec_4_T_3[5:0] ? myVec_40 : _GEN_3921; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3923 = 6'h29 == _myNewVec_4_T_3[5:0] ? myVec_41 : _GEN_3922; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3924 = 6'h2a == _myNewVec_4_T_3[5:0] ? myVec_42 : _GEN_3923; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3925 = 6'h2b == _myNewVec_4_T_3[5:0] ? myVec_43 : _GEN_3924; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3926 = 6'h2c == _myNewVec_4_T_3[5:0] ? myVec_44 : _GEN_3925; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3927 = 6'h2d == _myNewVec_4_T_3[5:0] ? myVec_45 : _GEN_3926; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3928 = 6'h2e == _myNewVec_4_T_3[5:0] ? myVec_46 : _GEN_3927; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3929 = 6'h2f == _myNewVec_4_T_3[5:0] ? myVec_47 : _GEN_3928; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3930 = 6'h30 == _myNewVec_4_T_3[5:0] ? myVec_48 : _GEN_3929; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3931 = 6'h31 == _myNewVec_4_T_3[5:0] ? myVec_49 : _GEN_3930; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3932 = 6'h32 == _myNewVec_4_T_3[5:0] ? myVec_50 : _GEN_3931; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3933 = 6'h33 == _myNewVec_4_T_3[5:0] ? myVec_51 : _GEN_3932; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3934 = 6'h34 == _myNewVec_4_T_3[5:0] ? myVec_52 : _GEN_3933; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3935 = 6'h35 == _myNewVec_4_T_3[5:0] ? myVec_53 : _GEN_3934; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3936 = 6'h36 == _myNewVec_4_T_3[5:0] ? myVec_54 : _GEN_3935; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3937 = 6'h37 == _myNewVec_4_T_3[5:0] ? myVec_55 : _GEN_3936; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3938 = 6'h38 == _myNewVec_4_T_3[5:0] ? myVec_56 : _GEN_3937; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3939 = 6'h39 == _myNewVec_4_T_3[5:0] ? myVec_57 : _GEN_3938; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3940 = 6'h3a == _myNewVec_4_T_3[5:0] ? myVec_58 : _GEN_3939; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3941 = 6'h3b == _myNewVec_4_T_3[5:0] ? myVec_59 : _GEN_3940; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3942 = 6'h3c == _myNewVec_4_T_3[5:0] ? myVec_60 : _GEN_3941; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3943 = 6'h3d == _myNewVec_4_T_3[5:0] ? myVec_61 : _GEN_3942; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3944 = 6'h3e == _myNewVec_4_T_3[5:0] ? myVec_62 : _GEN_3943; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_4 = 6'h3f == _myNewVec_4_T_3[5:0] ? myVec_63 : _GEN_3944; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_3_T_3 = _myNewVec_63_T_1 + 16'h3c; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_3947 = 6'h1 == _myNewVec_3_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3948 = 6'h2 == _myNewVec_3_T_3[5:0] ? myVec_2 : _GEN_3947; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3949 = 6'h3 == _myNewVec_3_T_3[5:0] ? myVec_3 : _GEN_3948; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3950 = 6'h4 == _myNewVec_3_T_3[5:0] ? myVec_4 : _GEN_3949; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3951 = 6'h5 == _myNewVec_3_T_3[5:0] ? myVec_5 : _GEN_3950; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3952 = 6'h6 == _myNewVec_3_T_3[5:0] ? myVec_6 : _GEN_3951; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3953 = 6'h7 == _myNewVec_3_T_3[5:0] ? myVec_7 : _GEN_3952; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3954 = 6'h8 == _myNewVec_3_T_3[5:0] ? myVec_8 : _GEN_3953; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3955 = 6'h9 == _myNewVec_3_T_3[5:0] ? myVec_9 : _GEN_3954; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3956 = 6'ha == _myNewVec_3_T_3[5:0] ? myVec_10 : _GEN_3955; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3957 = 6'hb == _myNewVec_3_T_3[5:0] ? myVec_11 : _GEN_3956; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3958 = 6'hc == _myNewVec_3_T_3[5:0] ? myVec_12 : _GEN_3957; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3959 = 6'hd == _myNewVec_3_T_3[5:0] ? myVec_13 : _GEN_3958; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3960 = 6'he == _myNewVec_3_T_3[5:0] ? myVec_14 : _GEN_3959; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3961 = 6'hf == _myNewVec_3_T_3[5:0] ? myVec_15 : _GEN_3960; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3962 = 6'h10 == _myNewVec_3_T_3[5:0] ? myVec_16 : _GEN_3961; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3963 = 6'h11 == _myNewVec_3_T_3[5:0] ? myVec_17 : _GEN_3962; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3964 = 6'h12 == _myNewVec_3_T_3[5:0] ? myVec_18 : _GEN_3963; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3965 = 6'h13 == _myNewVec_3_T_3[5:0] ? myVec_19 : _GEN_3964; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3966 = 6'h14 == _myNewVec_3_T_3[5:0] ? myVec_20 : _GEN_3965; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3967 = 6'h15 == _myNewVec_3_T_3[5:0] ? myVec_21 : _GEN_3966; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3968 = 6'h16 == _myNewVec_3_T_3[5:0] ? myVec_22 : _GEN_3967; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3969 = 6'h17 == _myNewVec_3_T_3[5:0] ? myVec_23 : _GEN_3968; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3970 = 6'h18 == _myNewVec_3_T_3[5:0] ? myVec_24 : _GEN_3969; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3971 = 6'h19 == _myNewVec_3_T_3[5:0] ? myVec_25 : _GEN_3970; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3972 = 6'h1a == _myNewVec_3_T_3[5:0] ? myVec_26 : _GEN_3971; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3973 = 6'h1b == _myNewVec_3_T_3[5:0] ? myVec_27 : _GEN_3972; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3974 = 6'h1c == _myNewVec_3_T_3[5:0] ? myVec_28 : _GEN_3973; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3975 = 6'h1d == _myNewVec_3_T_3[5:0] ? myVec_29 : _GEN_3974; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3976 = 6'h1e == _myNewVec_3_T_3[5:0] ? myVec_30 : _GEN_3975; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3977 = 6'h1f == _myNewVec_3_T_3[5:0] ? myVec_31 : _GEN_3976; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3978 = 6'h20 == _myNewVec_3_T_3[5:0] ? myVec_32 : _GEN_3977; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3979 = 6'h21 == _myNewVec_3_T_3[5:0] ? myVec_33 : _GEN_3978; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3980 = 6'h22 == _myNewVec_3_T_3[5:0] ? myVec_34 : _GEN_3979; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3981 = 6'h23 == _myNewVec_3_T_3[5:0] ? myVec_35 : _GEN_3980; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3982 = 6'h24 == _myNewVec_3_T_3[5:0] ? myVec_36 : _GEN_3981; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3983 = 6'h25 == _myNewVec_3_T_3[5:0] ? myVec_37 : _GEN_3982; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3984 = 6'h26 == _myNewVec_3_T_3[5:0] ? myVec_38 : _GEN_3983; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3985 = 6'h27 == _myNewVec_3_T_3[5:0] ? myVec_39 : _GEN_3984; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3986 = 6'h28 == _myNewVec_3_T_3[5:0] ? myVec_40 : _GEN_3985; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3987 = 6'h29 == _myNewVec_3_T_3[5:0] ? myVec_41 : _GEN_3986; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3988 = 6'h2a == _myNewVec_3_T_3[5:0] ? myVec_42 : _GEN_3987; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3989 = 6'h2b == _myNewVec_3_T_3[5:0] ? myVec_43 : _GEN_3988; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3990 = 6'h2c == _myNewVec_3_T_3[5:0] ? myVec_44 : _GEN_3989; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3991 = 6'h2d == _myNewVec_3_T_3[5:0] ? myVec_45 : _GEN_3990; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3992 = 6'h2e == _myNewVec_3_T_3[5:0] ? myVec_46 : _GEN_3991; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3993 = 6'h2f == _myNewVec_3_T_3[5:0] ? myVec_47 : _GEN_3992; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3994 = 6'h30 == _myNewVec_3_T_3[5:0] ? myVec_48 : _GEN_3993; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3995 = 6'h31 == _myNewVec_3_T_3[5:0] ? myVec_49 : _GEN_3994; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3996 = 6'h32 == _myNewVec_3_T_3[5:0] ? myVec_50 : _GEN_3995; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3997 = 6'h33 == _myNewVec_3_T_3[5:0] ? myVec_51 : _GEN_3996; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3998 = 6'h34 == _myNewVec_3_T_3[5:0] ? myVec_52 : _GEN_3997; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_3999 = 6'h35 == _myNewVec_3_T_3[5:0] ? myVec_53 : _GEN_3998; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4000 = 6'h36 == _myNewVec_3_T_3[5:0] ? myVec_54 : _GEN_3999; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4001 = 6'h37 == _myNewVec_3_T_3[5:0] ? myVec_55 : _GEN_4000; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4002 = 6'h38 == _myNewVec_3_T_3[5:0] ? myVec_56 : _GEN_4001; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4003 = 6'h39 == _myNewVec_3_T_3[5:0] ? myVec_57 : _GEN_4002; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4004 = 6'h3a == _myNewVec_3_T_3[5:0] ? myVec_58 : _GEN_4003; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4005 = 6'h3b == _myNewVec_3_T_3[5:0] ? myVec_59 : _GEN_4004; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4006 = 6'h3c == _myNewVec_3_T_3[5:0] ? myVec_60 : _GEN_4005; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4007 = 6'h3d == _myNewVec_3_T_3[5:0] ? myVec_61 : _GEN_4006; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4008 = 6'h3e == _myNewVec_3_T_3[5:0] ? myVec_62 : _GEN_4007; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_3 = 6'h3f == _myNewVec_3_T_3[5:0] ? myVec_63 : _GEN_4008; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_2_T_3 = _myNewVec_63_T_1 + 16'h3d; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4011 = 6'h1 == _myNewVec_2_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4012 = 6'h2 == _myNewVec_2_T_3[5:0] ? myVec_2 : _GEN_4011; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4013 = 6'h3 == _myNewVec_2_T_3[5:0] ? myVec_3 : _GEN_4012; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4014 = 6'h4 == _myNewVec_2_T_3[5:0] ? myVec_4 : _GEN_4013; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4015 = 6'h5 == _myNewVec_2_T_3[5:0] ? myVec_5 : _GEN_4014; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4016 = 6'h6 == _myNewVec_2_T_3[5:0] ? myVec_6 : _GEN_4015; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4017 = 6'h7 == _myNewVec_2_T_3[5:0] ? myVec_7 : _GEN_4016; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4018 = 6'h8 == _myNewVec_2_T_3[5:0] ? myVec_8 : _GEN_4017; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4019 = 6'h9 == _myNewVec_2_T_3[5:0] ? myVec_9 : _GEN_4018; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4020 = 6'ha == _myNewVec_2_T_3[5:0] ? myVec_10 : _GEN_4019; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4021 = 6'hb == _myNewVec_2_T_3[5:0] ? myVec_11 : _GEN_4020; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4022 = 6'hc == _myNewVec_2_T_3[5:0] ? myVec_12 : _GEN_4021; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4023 = 6'hd == _myNewVec_2_T_3[5:0] ? myVec_13 : _GEN_4022; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4024 = 6'he == _myNewVec_2_T_3[5:0] ? myVec_14 : _GEN_4023; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4025 = 6'hf == _myNewVec_2_T_3[5:0] ? myVec_15 : _GEN_4024; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4026 = 6'h10 == _myNewVec_2_T_3[5:0] ? myVec_16 : _GEN_4025; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4027 = 6'h11 == _myNewVec_2_T_3[5:0] ? myVec_17 : _GEN_4026; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4028 = 6'h12 == _myNewVec_2_T_3[5:0] ? myVec_18 : _GEN_4027; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4029 = 6'h13 == _myNewVec_2_T_3[5:0] ? myVec_19 : _GEN_4028; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4030 = 6'h14 == _myNewVec_2_T_3[5:0] ? myVec_20 : _GEN_4029; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4031 = 6'h15 == _myNewVec_2_T_3[5:0] ? myVec_21 : _GEN_4030; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4032 = 6'h16 == _myNewVec_2_T_3[5:0] ? myVec_22 : _GEN_4031; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4033 = 6'h17 == _myNewVec_2_T_3[5:0] ? myVec_23 : _GEN_4032; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4034 = 6'h18 == _myNewVec_2_T_3[5:0] ? myVec_24 : _GEN_4033; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4035 = 6'h19 == _myNewVec_2_T_3[5:0] ? myVec_25 : _GEN_4034; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4036 = 6'h1a == _myNewVec_2_T_3[5:0] ? myVec_26 : _GEN_4035; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4037 = 6'h1b == _myNewVec_2_T_3[5:0] ? myVec_27 : _GEN_4036; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4038 = 6'h1c == _myNewVec_2_T_3[5:0] ? myVec_28 : _GEN_4037; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4039 = 6'h1d == _myNewVec_2_T_3[5:0] ? myVec_29 : _GEN_4038; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4040 = 6'h1e == _myNewVec_2_T_3[5:0] ? myVec_30 : _GEN_4039; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4041 = 6'h1f == _myNewVec_2_T_3[5:0] ? myVec_31 : _GEN_4040; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4042 = 6'h20 == _myNewVec_2_T_3[5:0] ? myVec_32 : _GEN_4041; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4043 = 6'h21 == _myNewVec_2_T_3[5:0] ? myVec_33 : _GEN_4042; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4044 = 6'h22 == _myNewVec_2_T_3[5:0] ? myVec_34 : _GEN_4043; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4045 = 6'h23 == _myNewVec_2_T_3[5:0] ? myVec_35 : _GEN_4044; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4046 = 6'h24 == _myNewVec_2_T_3[5:0] ? myVec_36 : _GEN_4045; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4047 = 6'h25 == _myNewVec_2_T_3[5:0] ? myVec_37 : _GEN_4046; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4048 = 6'h26 == _myNewVec_2_T_3[5:0] ? myVec_38 : _GEN_4047; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4049 = 6'h27 == _myNewVec_2_T_3[5:0] ? myVec_39 : _GEN_4048; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4050 = 6'h28 == _myNewVec_2_T_3[5:0] ? myVec_40 : _GEN_4049; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4051 = 6'h29 == _myNewVec_2_T_3[5:0] ? myVec_41 : _GEN_4050; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4052 = 6'h2a == _myNewVec_2_T_3[5:0] ? myVec_42 : _GEN_4051; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4053 = 6'h2b == _myNewVec_2_T_3[5:0] ? myVec_43 : _GEN_4052; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4054 = 6'h2c == _myNewVec_2_T_3[5:0] ? myVec_44 : _GEN_4053; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4055 = 6'h2d == _myNewVec_2_T_3[5:0] ? myVec_45 : _GEN_4054; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4056 = 6'h2e == _myNewVec_2_T_3[5:0] ? myVec_46 : _GEN_4055; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4057 = 6'h2f == _myNewVec_2_T_3[5:0] ? myVec_47 : _GEN_4056; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4058 = 6'h30 == _myNewVec_2_T_3[5:0] ? myVec_48 : _GEN_4057; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4059 = 6'h31 == _myNewVec_2_T_3[5:0] ? myVec_49 : _GEN_4058; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4060 = 6'h32 == _myNewVec_2_T_3[5:0] ? myVec_50 : _GEN_4059; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4061 = 6'h33 == _myNewVec_2_T_3[5:0] ? myVec_51 : _GEN_4060; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4062 = 6'h34 == _myNewVec_2_T_3[5:0] ? myVec_52 : _GEN_4061; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4063 = 6'h35 == _myNewVec_2_T_3[5:0] ? myVec_53 : _GEN_4062; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4064 = 6'h36 == _myNewVec_2_T_3[5:0] ? myVec_54 : _GEN_4063; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4065 = 6'h37 == _myNewVec_2_T_3[5:0] ? myVec_55 : _GEN_4064; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4066 = 6'h38 == _myNewVec_2_T_3[5:0] ? myVec_56 : _GEN_4065; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4067 = 6'h39 == _myNewVec_2_T_3[5:0] ? myVec_57 : _GEN_4066; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4068 = 6'h3a == _myNewVec_2_T_3[5:0] ? myVec_58 : _GEN_4067; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4069 = 6'h3b == _myNewVec_2_T_3[5:0] ? myVec_59 : _GEN_4068; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4070 = 6'h3c == _myNewVec_2_T_3[5:0] ? myVec_60 : _GEN_4069; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4071 = 6'h3d == _myNewVec_2_T_3[5:0] ? myVec_61 : _GEN_4070; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4072 = 6'h3e == _myNewVec_2_T_3[5:0] ? myVec_62 : _GEN_4071; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_2 = 6'h3f == _myNewVec_2_T_3[5:0] ? myVec_63 : _GEN_4072; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_1_T_3 = _myNewVec_63_T_1 + 16'h3e; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4075 = 6'h1 == _myNewVec_1_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4076 = 6'h2 == _myNewVec_1_T_3[5:0] ? myVec_2 : _GEN_4075; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4077 = 6'h3 == _myNewVec_1_T_3[5:0] ? myVec_3 : _GEN_4076; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4078 = 6'h4 == _myNewVec_1_T_3[5:0] ? myVec_4 : _GEN_4077; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4079 = 6'h5 == _myNewVec_1_T_3[5:0] ? myVec_5 : _GEN_4078; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4080 = 6'h6 == _myNewVec_1_T_3[5:0] ? myVec_6 : _GEN_4079; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4081 = 6'h7 == _myNewVec_1_T_3[5:0] ? myVec_7 : _GEN_4080; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4082 = 6'h8 == _myNewVec_1_T_3[5:0] ? myVec_8 : _GEN_4081; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4083 = 6'h9 == _myNewVec_1_T_3[5:0] ? myVec_9 : _GEN_4082; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4084 = 6'ha == _myNewVec_1_T_3[5:0] ? myVec_10 : _GEN_4083; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4085 = 6'hb == _myNewVec_1_T_3[5:0] ? myVec_11 : _GEN_4084; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4086 = 6'hc == _myNewVec_1_T_3[5:0] ? myVec_12 : _GEN_4085; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4087 = 6'hd == _myNewVec_1_T_3[5:0] ? myVec_13 : _GEN_4086; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4088 = 6'he == _myNewVec_1_T_3[5:0] ? myVec_14 : _GEN_4087; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4089 = 6'hf == _myNewVec_1_T_3[5:0] ? myVec_15 : _GEN_4088; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4090 = 6'h10 == _myNewVec_1_T_3[5:0] ? myVec_16 : _GEN_4089; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4091 = 6'h11 == _myNewVec_1_T_3[5:0] ? myVec_17 : _GEN_4090; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4092 = 6'h12 == _myNewVec_1_T_3[5:0] ? myVec_18 : _GEN_4091; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4093 = 6'h13 == _myNewVec_1_T_3[5:0] ? myVec_19 : _GEN_4092; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4094 = 6'h14 == _myNewVec_1_T_3[5:0] ? myVec_20 : _GEN_4093; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4095 = 6'h15 == _myNewVec_1_T_3[5:0] ? myVec_21 : _GEN_4094; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4096 = 6'h16 == _myNewVec_1_T_3[5:0] ? myVec_22 : _GEN_4095; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4097 = 6'h17 == _myNewVec_1_T_3[5:0] ? myVec_23 : _GEN_4096; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4098 = 6'h18 == _myNewVec_1_T_3[5:0] ? myVec_24 : _GEN_4097; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4099 = 6'h19 == _myNewVec_1_T_3[5:0] ? myVec_25 : _GEN_4098; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4100 = 6'h1a == _myNewVec_1_T_3[5:0] ? myVec_26 : _GEN_4099; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4101 = 6'h1b == _myNewVec_1_T_3[5:0] ? myVec_27 : _GEN_4100; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4102 = 6'h1c == _myNewVec_1_T_3[5:0] ? myVec_28 : _GEN_4101; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4103 = 6'h1d == _myNewVec_1_T_3[5:0] ? myVec_29 : _GEN_4102; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4104 = 6'h1e == _myNewVec_1_T_3[5:0] ? myVec_30 : _GEN_4103; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4105 = 6'h1f == _myNewVec_1_T_3[5:0] ? myVec_31 : _GEN_4104; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4106 = 6'h20 == _myNewVec_1_T_3[5:0] ? myVec_32 : _GEN_4105; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4107 = 6'h21 == _myNewVec_1_T_3[5:0] ? myVec_33 : _GEN_4106; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4108 = 6'h22 == _myNewVec_1_T_3[5:0] ? myVec_34 : _GEN_4107; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4109 = 6'h23 == _myNewVec_1_T_3[5:0] ? myVec_35 : _GEN_4108; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4110 = 6'h24 == _myNewVec_1_T_3[5:0] ? myVec_36 : _GEN_4109; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4111 = 6'h25 == _myNewVec_1_T_3[5:0] ? myVec_37 : _GEN_4110; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4112 = 6'h26 == _myNewVec_1_T_3[5:0] ? myVec_38 : _GEN_4111; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4113 = 6'h27 == _myNewVec_1_T_3[5:0] ? myVec_39 : _GEN_4112; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4114 = 6'h28 == _myNewVec_1_T_3[5:0] ? myVec_40 : _GEN_4113; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4115 = 6'h29 == _myNewVec_1_T_3[5:0] ? myVec_41 : _GEN_4114; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4116 = 6'h2a == _myNewVec_1_T_3[5:0] ? myVec_42 : _GEN_4115; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4117 = 6'h2b == _myNewVec_1_T_3[5:0] ? myVec_43 : _GEN_4116; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4118 = 6'h2c == _myNewVec_1_T_3[5:0] ? myVec_44 : _GEN_4117; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4119 = 6'h2d == _myNewVec_1_T_3[5:0] ? myVec_45 : _GEN_4118; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4120 = 6'h2e == _myNewVec_1_T_3[5:0] ? myVec_46 : _GEN_4119; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4121 = 6'h2f == _myNewVec_1_T_3[5:0] ? myVec_47 : _GEN_4120; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4122 = 6'h30 == _myNewVec_1_T_3[5:0] ? myVec_48 : _GEN_4121; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4123 = 6'h31 == _myNewVec_1_T_3[5:0] ? myVec_49 : _GEN_4122; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4124 = 6'h32 == _myNewVec_1_T_3[5:0] ? myVec_50 : _GEN_4123; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4125 = 6'h33 == _myNewVec_1_T_3[5:0] ? myVec_51 : _GEN_4124; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4126 = 6'h34 == _myNewVec_1_T_3[5:0] ? myVec_52 : _GEN_4125; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4127 = 6'h35 == _myNewVec_1_T_3[5:0] ? myVec_53 : _GEN_4126; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4128 = 6'h36 == _myNewVec_1_T_3[5:0] ? myVec_54 : _GEN_4127; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4129 = 6'h37 == _myNewVec_1_T_3[5:0] ? myVec_55 : _GEN_4128; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4130 = 6'h38 == _myNewVec_1_T_3[5:0] ? myVec_56 : _GEN_4129; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4131 = 6'h39 == _myNewVec_1_T_3[5:0] ? myVec_57 : _GEN_4130; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4132 = 6'h3a == _myNewVec_1_T_3[5:0] ? myVec_58 : _GEN_4131; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4133 = 6'h3b == _myNewVec_1_T_3[5:0] ? myVec_59 : _GEN_4132; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4134 = 6'h3c == _myNewVec_1_T_3[5:0] ? myVec_60 : _GEN_4133; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4135 = 6'h3d == _myNewVec_1_T_3[5:0] ? myVec_61 : _GEN_4134; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4136 = 6'h3e == _myNewVec_1_T_3[5:0] ? myVec_62 : _GEN_4135; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_1 = 6'h3f == _myNewVec_1_T_3[5:0] ? myVec_63 : _GEN_4136; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [15:0] _myNewVec_0_T_3 = _myNewVec_63_T_1 + 16'h3f; // @[hh_datapath_chisel.scala 234:60]
  wire [31:0] _GEN_4139 = 6'h1 == _myNewVec_0_T_3[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4140 = 6'h2 == _myNewVec_0_T_3[5:0] ? myVec_2 : _GEN_4139; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4141 = 6'h3 == _myNewVec_0_T_3[5:0] ? myVec_3 : _GEN_4140; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4142 = 6'h4 == _myNewVec_0_T_3[5:0] ? myVec_4 : _GEN_4141; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4143 = 6'h5 == _myNewVec_0_T_3[5:0] ? myVec_5 : _GEN_4142; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4144 = 6'h6 == _myNewVec_0_T_3[5:0] ? myVec_6 : _GEN_4143; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4145 = 6'h7 == _myNewVec_0_T_3[5:0] ? myVec_7 : _GEN_4144; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4146 = 6'h8 == _myNewVec_0_T_3[5:0] ? myVec_8 : _GEN_4145; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4147 = 6'h9 == _myNewVec_0_T_3[5:0] ? myVec_9 : _GEN_4146; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4148 = 6'ha == _myNewVec_0_T_3[5:0] ? myVec_10 : _GEN_4147; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4149 = 6'hb == _myNewVec_0_T_3[5:0] ? myVec_11 : _GEN_4148; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4150 = 6'hc == _myNewVec_0_T_3[5:0] ? myVec_12 : _GEN_4149; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4151 = 6'hd == _myNewVec_0_T_3[5:0] ? myVec_13 : _GEN_4150; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4152 = 6'he == _myNewVec_0_T_3[5:0] ? myVec_14 : _GEN_4151; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4153 = 6'hf == _myNewVec_0_T_3[5:0] ? myVec_15 : _GEN_4152; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4154 = 6'h10 == _myNewVec_0_T_3[5:0] ? myVec_16 : _GEN_4153; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4155 = 6'h11 == _myNewVec_0_T_3[5:0] ? myVec_17 : _GEN_4154; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4156 = 6'h12 == _myNewVec_0_T_3[5:0] ? myVec_18 : _GEN_4155; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4157 = 6'h13 == _myNewVec_0_T_3[5:0] ? myVec_19 : _GEN_4156; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4158 = 6'h14 == _myNewVec_0_T_3[5:0] ? myVec_20 : _GEN_4157; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4159 = 6'h15 == _myNewVec_0_T_3[5:0] ? myVec_21 : _GEN_4158; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4160 = 6'h16 == _myNewVec_0_T_3[5:0] ? myVec_22 : _GEN_4159; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4161 = 6'h17 == _myNewVec_0_T_3[5:0] ? myVec_23 : _GEN_4160; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4162 = 6'h18 == _myNewVec_0_T_3[5:0] ? myVec_24 : _GEN_4161; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4163 = 6'h19 == _myNewVec_0_T_3[5:0] ? myVec_25 : _GEN_4162; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4164 = 6'h1a == _myNewVec_0_T_3[5:0] ? myVec_26 : _GEN_4163; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4165 = 6'h1b == _myNewVec_0_T_3[5:0] ? myVec_27 : _GEN_4164; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4166 = 6'h1c == _myNewVec_0_T_3[5:0] ? myVec_28 : _GEN_4165; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4167 = 6'h1d == _myNewVec_0_T_3[5:0] ? myVec_29 : _GEN_4166; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4168 = 6'h1e == _myNewVec_0_T_3[5:0] ? myVec_30 : _GEN_4167; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4169 = 6'h1f == _myNewVec_0_T_3[5:0] ? myVec_31 : _GEN_4168; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4170 = 6'h20 == _myNewVec_0_T_3[5:0] ? myVec_32 : _GEN_4169; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4171 = 6'h21 == _myNewVec_0_T_3[5:0] ? myVec_33 : _GEN_4170; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4172 = 6'h22 == _myNewVec_0_T_3[5:0] ? myVec_34 : _GEN_4171; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4173 = 6'h23 == _myNewVec_0_T_3[5:0] ? myVec_35 : _GEN_4172; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4174 = 6'h24 == _myNewVec_0_T_3[5:0] ? myVec_36 : _GEN_4173; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4175 = 6'h25 == _myNewVec_0_T_3[5:0] ? myVec_37 : _GEN_4174; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4176 = 6'h26 == _myNewVec_0_T_3[5:0] ? myVec_38 : _GEN_4175; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4177 = 6'h27 == _myNewVec_0_T_3[5:0] ? myVec_39 : _GEN_4176; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4178 = 6'h28 == _myNewVec_0_T_3[5:0] ? myVec_40 : _GEN_4177; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4179 = 6'h29 == _myNewVec_0_T_3[5:0] ? myVec_41 : _GEN_4178; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4180 = 6'h2a == _myNewVec_0_T_3[5:0] ? myVec_42 : _GEN_4179; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4181 = 6'h2b == _myNewVec_0_T_3[5:0] ? myVec_43 : _GEN_4180; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4182 = 6'h2c == _myNewVec_0_T_3[5:0] ? myVec_44 : _GEN_4181; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4183 = 6'h2d == _myNewVec_0_T_3[5:0] ? myVec_45 : _GEN_4182; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4184 = 6'h2e == _myNewVec_0_T_3[5:0] ? myVec_46 : _GEN_4183; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4185 = 6'h2f == _myNewVec_0_T_3[5:0] ? myVec_47 : _GEN_4184; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4186 = 6'h30 == _myNewVec_0_T_3[5:0] ? myVec_48 : _GEN_4185; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4187 = 6'h31 == _myNewVec_0_T_3[5:0] ? myVec_49 : _GEN_4186; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4188 = 6'h32 == _myNewVec_0_T_3[5:0] ? myVec_50 : _GEN_4187; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4189 = 6'h33 == _myNewVec_0_T_3[5:0] ? myVec_51 : _GEN_4188; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4190 = 6'h34 == _myNewVec_0_T_3[5:0] ? myVec_52 : _GEN_4189; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4191 = 6'h35 == _myNewVec_0_T_3[5:0] ? myVec_53 : _GEN_4190; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4192 = 6'h36 == _myNewVec_0_T_3[5:0] ? myVec_54 : _GEN_4191; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4193 = 6'h37 == _myNewVec_0_T_3[5:0] ? myVec_55 : _GEN_4192; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4194 = 6'h38 == _myNewVec_0_T_3[5:0] ? myVec_56 : _GEN_4193; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4195 = 6'h39 == _myNewVec_0_T_3[5:0] ? myVec_57 : _GEN_4194; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4196 = 6'h3a == _myNewVec_0_T_3[5:0] ? myVec_58 : _GEN_4195; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4197 = 6'h3b == _myNewVec_0_T_3[5:0] ? myVec_59 : _GEN_4196; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4198 = 6'h3c == _myNewVec_0_T_3[5:0] ? myVec_60 : _GEN_4197; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4199 = 6'h3d == _myNewVec_0_T_3[5:0] ? myVec_61 : _GEN_4198; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] _GEN_4200 = 6'h3e == _myNewVec_0_T_3[5:0] ? myVec_62 : _GEN_4199; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [31:0] myNewVec_0 = 6'h3f == _myNewVec_0_T_3[5:0] ? myVec_63 : _GEN_4200; // @[hh_datapath_chisel.scala 234:{37,37}]
  wire [255:0] myNewWire_lo_lo_lo = {myNewVec_7,myNewVec_6,myNewVec_5,myNewVec_4,myNewVec_3,myNewVec_2,myNewVec_1,
    myNewVec_0}; // @[hh_datapath_chisel.scala 238:27]
  wire [511:0] myNewWire_lo_lo = {myNewVec_15,myNewVec_14,myNewVec_13,myNewVec_12,myNewVec_11,myNewVec_10,myNewVec_9,
    myNewVec_8,myNewWire_lo_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [1023:0] myNewWire_lo = {myNewVec_31,myNewVec_30,myNewVec_29,myNewVec_28,myNewVec_27,myNewVec_26,myNewVec_25,
    myNewVec_24,myNewWire_lo_hi_lo,myNewWire_lo_lo}; // @[hh_datapath_chisel.scala 238:27]
  wire [2079:0] _vk_update_T = {vk1,myNewWire_hi,myNewWire_lo}; // @[Cat.scala 31:58]
  wire [21:0] _vk_update_T_3 = _myNewVec_63_T_1 * 6'h20; // @[hh_datapath_chisel.scala 242:57]
  wire [2079:0] _vk_update_T_4 = _vk_update_T >> _vk_update_T_3; // @[hh_datapath_chisel.scala 242:39]
  wire [2079:0] _GEN_4202 = io_vk1_vld ? _vk_update_T_4 : 2080'h0; // @[hh_datapath_chisel.scala 241:27 242:17 245:17]
  wire [2079:0] _GEN_4203 = io_rst ? 2080'h0 : _GEN_4202; // @[hh_datapath_chisel.scala 239:17 240:17]
  wire [2047:0] vk_update = _GEN_4203[2047:0]; // @[hh_datapath_chisel.scala 81:25]
  wire [2047:0] vk = io_vk1_vld ? vk_update : vk_reg; // @[hh_datapath_chisel.scala 155:21 156:10 158:10]
  wire [31:0] ddot_dout = FP_DDOT_dp_io_out_s; // @[hh_datapath_chisel.scala 254:15 75:25]
  wire [31:0] _GEN_41 = 6'h1 == io_hh_cnt[5:0] ? myVec_1 : myVec_0; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_42 = 6'h2 == io_hh_cnt[5:0] ? myVec_2 : _GEN_41; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_43 = 6'h3 == io_hh_cnt[5:0] ? myVec_3 : _GEN_42; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_44 = 6'h4 == io_hh_cnt[5:0] ? myVec_4 : _GEN_43; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_45 = 6'h5 == io_hh_cnt[5:0] ? myVec_5 : _GEN_44; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_46 = 6'h6 == io_hh_cnt[5:0] ? myVec_6 : _GEN_45; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_47 = 6'h7 == io_hh_cnt[5:0] ? myVec_7 : _GEN_46; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_48 = 6'h8 == io_hh_cnt[5:0] ? myVec_8 : _GEN_47; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_49 = 6'h9 == io_hh_cnt[5:0] ? myVec_9 : _GEN_48; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_50 = 6'ha == io_hh_cnt[5:0] ? myVec_10 : _GEN_49; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_51 = 6'hb == io_hh_cnt[5:0] ? myVec_11 : _GEN_50; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_52 = 6'hc == io_hh_cnt[5:0] ? myVec_12 : _GEN_51; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_53 = 6'hd == io_hh_cnt[5:0] ? myVec_13 : _GEN_52; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_54 = 6'he == io_hh_cnt[5:0] ? myVec_14 : _GEN_53; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_55 = 6'hf == io_hh_cnt[5:0] ? myVec_15 : _GEN_54; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_56 = 6'h10 == io_hh_cnt[5:0] ? myVec_16 : _GEN_55; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_57 = 6'h11 == io_hh_cnt[5:0] ? myVec_17 : _GEN_56; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_58 = 6'h12 == io_hh_cnt[5:0] ? myVec_18 : _GEN_57; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_59 = 6'h13 == io_hh_cnt[5:0] ? myVec_19 : _GEN_58; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_60 = 6'h14 == io_hh_cnt[5:0] ? myVec_20 : _GEN_59; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_61 = 6'h15 == io_hh_cnt[5:0] ? myVec_21 : _GEN_60; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_62 = 6'h16 == io_hh_cnt[5:0] ? myVec_22 : _GEN_61; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_63 = 6'h17 == io_hh_cnt[5:0] ? myVec_23 : _GEN_62; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_64 = 6'h18 == io_hh_cnt[5:0] ? myVec_24 : _GEN_63; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_65 = 6'h19 == io_hh_cnt[5:0] ? myVec_25 : _GEN_64; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_66 = 6'h1a == io_hh_cnt[5:0] ? myVec_26 : _GEN_65; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_67 = 6'h1b == io_hh_cnt[5:0] ? myVec_27 : _GEN_66; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_68 = 6'h1c == io_hh_cnt[5:0] ? myVec_28 : _GEN_67; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_69 = 6'h1d == io_hh_cnt[5:0] ? myVec_29 : _GEN_68; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_70 = 6'h1e == io_hh_cnt[5:0] ? myVec_30 : _GEN_69; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_71 = 6'h1f == io_hh_cnt[5:0] ? myVec_31 : _GEN_70; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_72 = 6'h20 == io_hh_cnt[5:0] ? myVec_32 : _GEN_71; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_73 = 6'h21 == io_hh_cnt[5:0] ? myVec_33 : _GEN_72; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_74 = 6'h22 == io_hh_cnt[5:0] ? myVec_34 : _GEN_73; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_75 = 6'h23 == io_hh_cnt[5:0] ? myVec_35 : _GEN_74; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_76 = 6'h24 == io_hh_cnt[5:0] ? myVec_36 : _GEN_75; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_77 = 6'h25 == io_hh_cnt[5:0] ? myVec_37 : _GEN_76; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_78 = 6'h26 == io_hh_cnt[5:0] ? myVec_38 : _GEN_77; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_79 = 6'h27 == io_hh_cnt[5:0] ? myVec_39 : _GEN_78; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_80 = 6'h28 == io_hh_cnt[5:0] ? myVec_40 : _GEN_79; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_81 = 6'h29 == io_hh_cnt[5:0] ? myVec_41 : _GEN_80; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_82 = 6'h2a == io_hh_cnt[5:0] ? myVec_42 : _GEN_81; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_83 = 6'h2b == io_hh_cnt[5:0] ? myVec_43 : _GEN_82; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_84 = 6'h2c == io_hh_cnt[5:0] ? myVec_44 : _GEN_83; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_85 = 6'h2d == io_hh_cnt[5:0] ? myVec_45 : _GEN_84; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_86 = 6'h2e == io_hh_cnt[5:0] ? myVec_46 : _GEN_85; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_87 = 6'h2f == io_hh_cnt[5:0] ? myVec_47 : _GEN_86; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_88 = 6'h30 == io_hh_cnt[5:0] ? myVec_48 : _GEN_87; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_89 = 6'h31 == io_hh_cnt[5:0] ? myVec_49 : _GEN_88; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_90 = 6'h32 == io_hh_cnt[5:0] ? myVec_50 : _GEN_89; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_91 = 6'h33 == io_hh_cnt[5:0] ? myVec_51 : _GEN_90; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_92 = 6'h34 == io_hh_cnt[5:0] ? myVec_52 : _GEN_91; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_93 = 6'h35 == io_hh_cnt[5:0] ? myVec_53 : _GEN_92; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_94 = 6'h36 == io_hh_cnt[5:0] ? myVec_54 : _GEN_93; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_95 = 6'h37 == io_hh_cnt[5:0] ? myVec_55 : _GEN_94; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_96 = 6'h38 == io_hh_cnt[5:0] ? myVec_56 : _GEN_95; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_97 = 6'h39 == io_hh_cnt[5:0] ? myVec_57 : _GEN_96; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_98 = 6'h3a == io_hh_cnt[5:0] ? myVec_58 : _GEN_97; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_99 = 6'h3b == io_hh_cnt[5:0] ? myVec_59 : _GEN_98; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_100 = 6'h3c == io_hh_cnt[5:0] ? myVec_60 : _GEN_99; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_101 = 6'h3d == io_hh_cnt[5:0] ? myVec_61 : _GEN_100; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_102 = 6'h3e == io_hh_cnt[5:0] ? myVec_62 : _GEN_101; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_103 = 6'h3f == io_hh_cnt[5:0] ? myVec_63 : _GEN_102; // @[hh_datapath_chisel.scala 226:{17,17}]
  wire [31:0] _GEN_104 = io_d1_rdy ? _GEN_103 : 32'h0; // @[hh_datapath_chisel.scala 225:26 226:17 228:17]
  wire [31:0] x1_update = io_rst ? 32'h0 : _GEN_104; // @[hh_datapath_chisel.scala 223:17 224:17]
  wire [31:0] d2_update = FP_square_root_newfpu_io_out_s; // @[hh_datapath_chisel.scala 259:15 90:25]
  wire [31:0] tk_update = hqr7_io_out_s; // @[hh_datapath_chisel.scala 268:14 92:25]
  wire [31:0] d5_update = FP_multiplier_10ccs_io_out_s; // @[hh_datapath_chisel.scala 274:14 94:25]
  reg [4063:0] d4_update_reg; // @[hh_datapath_chisel.scala 161:28]
  wire [4095:0] _d4_update_reg_T = {ddot_dout,d4_update_reg}; // @[Cat.scala 31:58]
  reg [31:0] myAxpyVec_0; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_1; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_2; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_3; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_4; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_5; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_6; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_7; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_8; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_9; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_10; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_11; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_12; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_13; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_14; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_15; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_16; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_17; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_18; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_19; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_20; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_21; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_22; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_23; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_24; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_25; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_26; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_27; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_28; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_29; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_30; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_31; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_32; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_33; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_34; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_35; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_36; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_37; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_38; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_39; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_40; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_41; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_42; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_43; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_44; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_45; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_46; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_47; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_48; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_49; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_50; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_51; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_52; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_53; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_54; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_55; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_56; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_57; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_58; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_59; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_60; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_61; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_62; // @[hh_datapath_chisel.scala 282:23]
  reg [31:0] myAxpyVec_63; // @[hh_datapath_chisel.scala 282:23]
  wire [255:0] io_hh_dout_lo_lo_lo = {myAxpyVec_7,myAxpyVec_6,myAxpyVec_5,myAxpyVec_4,myAxpyVec_3,myAxpyVec_2,
    myAxpyVec_1,myAxpyVec_0}; // @[hh_datapath_chisel.scala 290:28]
  wire [511:0] io_hh_dout_lo_lo = {myAxpyVec_15,myAxpyVec_14,myAxpyVec_13,myAxpyVec_12,myAxpyVec_11,myAxpyVec_10,
    myAxpyVec_9,myAxpyVec_8,io_hh_dout_lo_lo_lo}; // @[hh_datapath_chisel.scala 290:28]
  wire [255:0] io_hh_dout_lo_hi_lo = {myAxpyVec_23,myAxpyVec_22,myAxpyVec_21,myAxpyVec_20,myAxpyVec_19,myAxpyVec_18,
    myAxpyVec_17,myAxpyVec_16}; // @[hh_datapath_chisel.scala 290:28]
  wire [1023:0] io_hh_dout_lo = {myAxpyVec_31,myAxpyVec_30,myAxpyVec_29,myAxpyVec_28,myAxpyVec_27,myAxpyVec_26,
    myAxpyVec_25,myAxpyVec_24,io_hh_dout_lo_hi_lo,io_hh_dout_lo_lo}; // @[hh_datapath_chisel.scala 290:28]
  wire [255:0] io_hh_dout_hi_lo_lo = {myAxpyVec_39,myAxpyVec_38,myAxpyVec_37,myAxpyVec_36,myAxpyVec_35,myAxpyVec_34,
    myAxpyVec_33,myAxpyVec_32}; // @[hh_datapath_chisel.scala 290:28]
  wire [511:0] io_hh_dout_hi_lo = {myAxpyVec_47,myAxpyVec_46,myAxpyVec_45,myAxpyVec_44,myAxpyVec_43,myAxpyVec_42,
    myAxpyVec_41,myAxpyVec_40,io_hh_dout_hi_lo_lo}; // @[hh_datapath_chisel.scala 290:28]
  wire [255:0] io_hh_dout_hi_hi_lo = {myAxpyVec_55,myAxpyVec_54,myAxpyVec_53,myAxpyVec_52,myAxpyVec_51,myAxpyVec_50,
    myAxpyVec_49,myAxpyVec_48}; // @[hh_datapath_chisel.scala 290:28]
  wire [1023:0] io_hh_dout_hi = {myAxpyVec_63,myAxpyVec_62,myAxpyVec_61,myAxpyVec_60,myAxpyVec_59,myAxpyVec_58,
    myAxpyVec_57,myAxpyVec_56,io_hh_dout_hi_hi_lo,io_hh_dout_hi_lo}; // @[hh_datapath_chisel.scala 290:28]
  FP_DDOT_dp FP_DDOT_dp ( // @[hh_datapath_chisel.scala 248:21]
    .clock(FP_DDOT_dp_clock),
    .reset(FP_DDOT_dp_reset),
    .io_in_a_0(FP_DDOT_dp_io_in_a_0),
    .io_in_a_1(FP_DDOT_dp_io_in_a_1),
    .io_in_a_2(FP_DDOT_dp_io_in_a_2),
    .io_in_a_3(FP_DDOT_dp_io_in_a_3),
    .io_in_a_4(FP_DDOT_dp_io_in_a_4),
    .io_in_a_5(FP_DDOT_dp_io_in_a_5),
    .io_in_a_6(FP_DDOT_dp_io_in_a_6),
    .io_in_a_7(FP_DDOT_dp_io_in_a_7),
    .io_in_a_8(FP_DDOT_dp_io_in_a_8),
    .io_in_a_9(FP_DDOT_dp_io_in_a_9),
    .io_in_a_10(FP_DDOT_dp_io_in_a_10),
    .io_in_a_11(FP_DDOT_dp_io_in_a_11),
    .io_in_a_12(FP_DDOT_dp_io_in_a_12),
    .io_in_a_13(FP_DDOT_dp_io_in_a_13),
    .io_in_a_14(FP_DDOT_dp_io_in_a_14),
    .io_in_a_15(FP_DDOT_dp_io_in_a_15),
    .io_in_a_16(FP_DDOT_dp_io_in_a_16),
    .io_in_a_17(FP_DDOT_dp_io_in_a_17),
    .io_in_a_18(FP_DDOT_dp_io_in_a_18),
    .io_in_a_19(FP_DDOT_dp_io_in_a_19),
    .io_in_a_20(FP_DDOT_dp_io_in_a_20),
    .io_in_a_21(FP_DDOT_dp_io_in_a_21),
    .io_in_a_22(FP_DDOT_dp_io_in_a_22),
    .io_in_a_23(FP_DDOT_dp_io_in_a_23),
    .io_in_a_24(FP_DDOT_dp_io_in_a_24),
    .io_in_a_25(FP_DDOT_dp_io_in_a_25),
    .io_in_a_26(FP_DDOT_dp_io_in_a_26),
    .io_in_a_27(FP_DDOT_dp_io_in_a_27),
    .io_in_a_28(FP_DDOT_dp_io_in_a_28),
    .io_in_a_29(FP_DDOT_dp_io_in_a_29),
    .io_in_a_30(FP_DDOT_dp_io_in_a_30),
    .io_in_a_31(FP_DDOT_dp_io_in_a_31),
    .io_in_a_32(FP_DDOT_dp_io_in_a_32),
    .io_in_a_33(FP_DDOT_dp_io_in_a_33),
    .io_in_a_34(FP_DDOT_dp_io_in_a_34),
    .io_in_a_35(FP_DDOT_dp_io_in_a_35),
    .io_in_a_36(FP_DDOT_dp_io_in_a_36),
    .io_in_a_37(FP_DDOT_dp_io_in_a_37),
    .io_in_a_38(FP_DDOT_dp_io_in_a_38),
    .io_in_a_39(FP_DDOT_dp_io_in_a_39),
    .io_in_a_40(FP_DDOT_dp_io_in_a_40),
    .io_in_a_41(FP_DDOT_dp_io_in_a_41),
    .io_in_a_42(FP_DDOT_dp_io_in_a_42),
    .io_in_a_43(FP_DDOT_dp_io_in_a_43),
    .io_in_a_44(FP_DDOT_dp_io_in_a_44),
    .io_in_a_45(FP_DDOT_dp_io_in_a_45),
    .io_in_a_46(FP_DDOT_dp_io_in_a_46),
    .io_in_a_47(FP_DDOT_dp_io_in_a_47),
    .io_in_a_48(FP_DDOT_dp_io_in_a_48),
    .io_in_a_49(FP_DDOT_dp_io_in_a_49),
    .io_in_a_50(FP_DDOT_dp_io_in_a_50),
    .io_in_a_51(FP_DDOT_dp_io_in_a_51),
    .io_in_a_52(FP_DDOT_dp_io_in_a_52),
    .io_in_a_53(FP_DDOT_dp_io_in_a_53),
    .io_in_a_54(FP_DDOT_dp_io_in_a_54),
    .io_in_a_55(FP_DDOT_dp_io_in_a_55),
    .io_in_a_56(FP_DDOT_dp_io_in_a_56),
    .io_in_a_57(FP_DDOT_dp_io_in_a_57),
    .io_in_a_58(FP_DDOT_dp_io_in_a_58),
    .io_in_a_59(FP_DDOT_dp_io_in_a_59),
    .io_in_a_60(FP_DDOT_dp_io_in_a_60),
    .io_in_a_61(FP_DDOT_dp_io_in_a_61),
    .io_in_a_62(FP_DDOT_dp_io_in_a_62),
    .io_in_a_63(FP_DDOT_dp_io_in_a_63),
    .io_in_b_0(FP_DDOT_dp_io_in_b_0),
    .io_in_b_1(FP_DDOT_dp_io_in_b_1),
    .io_in_b_2(FP_DDOT_dp_io_in_b_2),
    .io_in_b_3(FP_DDOT_dp_io_in_b_3),
    .io_in_b_4(FP_DDOT_dp_io_in_b_4),
    .io_in_b_5(FP_DDOT_dp_io_in_b_5),
    .io_in_b_6(FP_DDOT_dp_io_in_b_6),
    .io_in_b_7(FP_DDOT_dp_io_in_b_7),
    .io_in_b_8(FP_DDOT_dp_io_in_b_8),
    .io_in_b_9(FP_DDOT_dp_io_in_b_9),
    .io_in_b_10(FP_DDOT_dp_io_in_b_10),
    .io_in_b_11(FP_DDOT_dp_io_in_b_11),
    .io_in_b_12(FP_DDOT_dp_io_in_b_12),
    .io_in_b_13(FP_DDOT_dp_io_in_b_13),
    .io_in_b_14(FP_DDOT_dp_io_in_b_14),
    .io_in_b_15(FP_DDOT_dp_io_in_b_15),
    .io_in_b_16(FP_DDOT_dp_io_in_b_16),
    .io_in_b_17(FP_DDOT_dp_io_in_b_17),
    .io_in_b_18(FP_DDOT_dp_io_in_b_18),
    .io_in_b_19(FP_DDOT_dp_io_in_b_19),
    .io_in_b_20(FP_DDOT_dp_io_in_b_20),
    .io_in_b_21(FP_DDOT_dp_io_in_b_21),
    .io_in_b_22(FP_DDOT_dp_io_in_b_22),
    .io_in_b_23(FP_DDOT_dp_io_in_b_23),
    .io_in_b_24(FP_DDOT_dp_io_in_b_24),
    .io_in_b_25(FP_DDOT_dp_io_in_b_25),
    .io_in_b_26(FP_DDOT_dp_io_in_b_26),
    .io_in_b_27(FP_DDOT_dp_io_in_b_27),
    .io_in_b_28(FP_DDOT_dp_io_in_b_28),
    .io_in_b_29(FP_DDOT_dp_io_in_b_29),
    .io_in_b_30(FP_DDOT_dp_io_in_b_30),
    .io_in_b_31(FP_DDOT_dp_io_in_b_31),
    .io_in_b_32(FP_DDOT_dp_io_in_b_32),
    .io_in_b_33(FP_DDOT_dp_io_in_b_33),
    .io_in_b_34(FP_DDOT_dp_io_in_b_34),
    .io_in_b_35(FP_DDOT_dp_io_in_b_35),
    .io_in_b_36(FP_DDOT_dp_io_in_b_36),
    .io_in_b_37(FP_DDOT_dp_io_in_b_37),
    .io_in_b_38(FP_DDOT_dp_io_in_b_38),
    .io_in_b_39(FP_DDOT_dp_io_in_b_39),
    .io_in_b_40(FP_DDOT_dp_io_in_b_40),
    .io_in_b_41(FP_DDOT_dp_io_in_b_41),
    .io_in_b_42(FP_DDOT_dp_io_in_b_42),
    .io_in_b_43(FP_DDOT_dp_io_in_b_43),
    .io_in_b_44(FP_DDOT_dp_io_in_b_44),
    .io_in_b_45(FP_DDOT_dp_io_in_b_45),
    .io_in_b_46(FP_DDOT_dp_io_in_b_46),
    .io_in_b_47(FP_DDOT_dp_io_in_b_47),
    .io_in_b_48(FP_DDOT_dp_io_in_b_48),
    .io_in_b_49(FP_DDOT_dp_io_in_b_49),
    .io_in_b_50(FP_DDOT_dp_io_in_b_50),
    .io_in_b_51(FP_DDOT_dp_io_in_b_51),
    .io_in_b_52(FP_DDOT_dp_io_in_b_52),
    .io_in_b_53(FP_DDOT_dp_io_in_b_53),
    .io_in_b_54(FP_DDOT_dp_io_in_b_54),
    .io_in_b_55(FP_DDOT_dp_io_in_b_55),
    .io_in_b_56(FP_DDOT_dp_io_in_b_56),
    .io_in_b_57(FP_DDOT_dp_io_in_b_57),
    .io_in_b_58(FP_DDOT_dp_io_in_b_58),
    .io_in_b_59(FP_DDOT_dp_io_in_b_59),
    .io_in_b_60(FP_DDOT_dp_io_in_b_60),
    .io_in_b_61(FP_DDOT_dp_io_in_b_61),
    .io_in_b_62(FP_DDOT_dp_io_in_b_62),
    .io_in_b_63(FP_DDOT_dp_io_in_b_63),
    .io_out_s(FP_DDOT_dp_io_out_s)
  );
  FP_square_root_newfpu FP_square_root_newfpu ( // @[hh_datapath_chisel.scala 256:22]
    .clock(FP_square_root_newfpu_clock),
    .reset(FP_square_root_newfpu_reset),
    .io_in_a(FP_square_root_newfpu_io_in_a),
    .io_out_s(FP_square_root_newfpu_io_out_s)
  );
  hqr5 hqr5 ( // @[hh_datapath_chisel.scala 261:20]
    .clock(hqr5_clock),
    .reset(hqr5_reset),
    .io_in_a(hqr5_io_in_a),
    .io_in_b(hqr5_io_in_b),
    .io_out_s(hqr5_io_out_s)
  );
  hqr7 hqr7 ( // @[hh_datapath_chisel.scala 266:20]
    .clock(hqr7_clock),
    .reset(hqr7_reset),
    .io_in_a(hqr7_io_in_a),
    .io_out_s(hqr7_io_out_s)
  );
  FP_multiplier_10ccs FP_multiplier_10ccs ( // @[hh_datapath_chisel.scala 270:21]
    .clock(FP_multiplier_10ccs_clock),
    .reset(FP_multiplier_10ccs_reset),
    .io_in_a(FP_multiplier_10ccs_io_in_a),
    .io_in_b(FP_multiplier_10ccs_io_in_b),
    .io_out_s(FP_multiplier_10ccs_io_out_s)
  );
  axpy_dp axpy_dp ( // @[hh_datapath_chisel.scala 276:20]
    .clock(axpy_dp_clock),
    .reset(axpy_dp_reset),
    .io_in_a(axpy_dp_io_in_a),
    .io_in_b_0(axpy_dp_io_in_b_0),
    .io_in_b_1(axpy_dp_io_in_b_1),
    .io_in_b_2(axpy_dp_io_in_b_2),
    .io_in_b_3(axpy_dp_io_in_b_3),
    .io_in_b_4(axpy_dp_io_in_b_4),
    .io_in_b_5(axpy_dp_io_in_b_5),
    .io_in_b_6(axpy_dp_io_in_b_6),
    .io_in_b_7(axpy_dp_io_in_b_7),
    .io_in_b_8(axpy_dp_io_in_b_8),
    .io_in_b_9(axpy_dp_io_in_b_9),
    .io_in_b_10(axpy_dp_io_in_b_10),
    .io_in_b_11(axpy_dp_io_in_b_11),
    .io_in_b_12(axpy_dp_io_in_b_12),
    .io_in_b_13(axpy_dp_io_in_b_13),
    .io_in_b_14(axpy_dp_io_in_b_14),
    .io_in_b_15(axpy_dp_io_in_b_15),
    .io_in_b_16(axpy_dp_io_in_b_16),
    .io_in_b_17(axpy_dp_io_in_b_17),
    .io_in_b_18(axpy_dp_io_in_b_18),
    .io_in_b_19(axpy_dp_io_in_b_19),
    .io_in_b_20(axpy_dp_io_in_b_20),
    .io_in_b_21(axpy_dp_io_in_b_21),
    .io_in_b_22(axpy_dp_io_in_b_22),
    .io_in_b_23(axpy_dp_io_in_b_23),
    .io_in_b_24(axpy_dp_io_in_b_24),
    .io_in_b_25(axpy_dp_io_in_b_25),
    .io_in_b_26(axpy_dp_io_in_b_26),
    .io_in_b_27(axpy_dp_io_in_b_27),
    .io_in_b_28(axpy_dp_io_in_b_28),
    .io_in_b_29(axpy_dp_io_in_b_29),
    .io_in_b_30(axpy_dp_io_in_b_30),
    .io_in_b_31(axpy_dp_io_in_b_31),
    .io_in_b_32(axpy_dp_io_in_b_32),
    .io_in_b_33(axpy_dp_io_in_b_33),
    .io_in_b_34(axpy_dp_io_in_b_34),
    .io_in_b_35(axpy_dp_io_in_b_35),
    .io_in_b_36(axpy_dp_io_in_b_36),
    .io_in_b_37(axpy_dp_io_in_b_37),
    .io_in_b_38(axpy_dp_io_in_b_38),
    .io_in_b_39(axpy_dp_io_in_b_39),
    .io_in_b_40(axpy_dp_io_in_b_40),
    .io_in_b_41(axpy_dp_io_in_b_41),
    .io_in_b_42(axpy_dp_io_in_b_42),
    .io_in_b_43(axpy_dp_io_in_b_43),
    .io_in_b_44(axpy_dp_io_in_b_44),
    .io_in_b_45(axpy_dp_io_in_b_45),
    .io_in_b_46(axpy_dp_io_in_b_46),
    .io_in_b_47(axpy_dp_io_in_b_47),
    .io_in_b_48(axpy_dp_io_in_b_48),
    .io_in_b_49(axpy_dp_io_in_b_49),
    .io_in_b_50(axpy_dp_io_in_b_50),
    .io_in_b_51(axpy_dp_io_in_b_51),
    .io_in_b_52(axpy_dp_io_in_b_52),
    .io_in_b_53(axpy_dp_io_in_b_53),
    .io_in_b_54(axpy_dp_io_in_b_54),
    .io_in_b_55(axpy_dp_io_in_b_55),
    .io_in_b_56(axpy_dp_io_in_b_56),
    .io_in_b_57(axpy_dp_io_in_b_57),
    .io_in_b_58(axpy_dp_io_in_b_58),
    .io_in_b_59(axpy_dp_io_in_b_59),
    .io_in_b_60(axpy_dp_io_in_b_60),
    .io_in_b_61(axpy_dp_io_in_b_61),
    .io_in_b_62(axpy_dp_io_in_b_62),
    .io_in_b_63(axpy_dp_io_in_b_63),
    .io_in_c_0(axpy_dp_io_in_c_0),
    .io_in_c_1(axpy_dp_io_in_c_1),
    .io_in_c_2(axpy_dp_io_in_c_2),
    .io_in_c_3(axpy_dp_io_in_c_3),
    .io_in_c_4(axpy_dp_io_in_c_4),
    .io_in_c_5(axpy_dp_io_in_c_5),
    .io_in_c_6(axpy_dp_io_in_c_6),
    .io_in_c_7(axpy_dp_io_in_c_7),
    .io_in_c_8(axpy_dp_io_in_c_8),
    .io_in_c_9(axpy_dp_io_in_c_9),
    .io_in_c_10(axpy_dp_io_in_c_10),
    .io_in_c_11(axpy_dp_io_in_c_11),
    .io_in_c_12(axpy_dp_io_in_c_12),
    .io_in_c_13(axpy_dp_io_in_c_13),
    .io_in_c_14(axpy_dp_io_in_c_14),
    .io_in_c_15(axpy_dp_io_in_c_15),
    .io_in_c_16(axpy_dp_io_in_c_16),
    .io_in_c_17(axpy_dp_io_in_c_17),
    .io_in_c_18(axpy_dp_io_in_c_18),
    .io_in_c_19(axpy_dp_io_in_c_19),
    .io_in_c_20(axpy_dp_io_in_c_20),
    .io_in_c_21(axpy_dp_io_in_c_21),
    .io_in_c_22(axpy_dp_io_in_c_22),
    .io_in_c_23(axpy_dp_io_in_c_23),
    .io_in_c_24(axpy_dp_io_in_c_24),
    .io_in_c_25(axpy_dp_io_in_c_25),
    .io_in_c_26(axpy_dp_io_in_c_26),
    .io_in_c_27(axpy_dp_io_in_c_27),
    .io_in_c_28(axpy_dp_io_in_c_28),
    .io_in_c_29(axpy_dp_io_in_c_29),
    .io_in_c_30(axpy_dp_io_in_c_30),
    .io_in_c_31(axpy_dp_io_in_c_31),
    .io_in_c_32(axpy_dp_io_in_c_32),
    .io_in_c_33(axpy_dp_io_in_c_33),
    .io_in_c_34(axpy_dp_io_in_c_34),
    .io_in_c_35(axpy_dp_io_in_c_35),
    .io_in_c_36(axpy_dp_io_in_c_36),
    .io_in_c_37(axpy_dp_io_in_c_37),
    .io_in_c_38(axpy_dp_io_in_c_38),
    .io_in_c_39(axpy_dp_io_in_c_39),
    .io_in_c_40(axpy_dp_io_in_c_40),
    .io_in_c_41(axpy_dp_io_in_c_41),
    .io_in_c_42(axpy_dp_io_in_c_42),
    .io_in_c_43(axpy_dp_io_in_c_43),
    .io_in_c_44(axpy_dp_io_in_c_44),
    .io_in_c_45(axpy_dp_io_in_c_45),
    .io_in_c_46(axpy_dp_io_in_c_46),
    .io_in_c_47(axpy_dp_io_in_c_47),
    .io_in_c_48(axpy_dp_io_in_c_48),
    .io_in_c_49(axpy_dp_io_in_c_49),
    .io_in_c_50(axpy_dp_io_in_c_50),
    .io_in_c_51(axpy_dp_io_in_c_51),
    .io_in_c_52(axpy_dp_io_in_c_52),
    .io_in_c_53(axpy_dp_io_in_c_53),
    .io_in_c_54(axpy_dp_io_in_c_54),
    .io_in_c_55(axpy_dp_io_in_c_55),
    .io_in_c_56(axpy_dp_io_in_c_56),
    .io_in_c_57(axpy_dp_io_in_c_57),
    .io_in_c_58(axpy_dp_io_in_c_58),
    .io_in_c_59(axpy_dp_io_in_c_59),
    .io_in_c_60(axpy_dp_io_in_c_60),
    .io_in_c_61(axpy_dp_io_in_c_61),
    .io_in_c_62(axpy_dp_io_in_c_62),
    .io_in_c_63(axpy_dp_io_in_c_63),
    .io_out_s_0(axpy_dp_io_out_s_0),
    .io_out_s_1(axpy_dp_io_out_s_1),
    .io_out_s_2(axpy_dp_io_out_s_2),
    .io_out_s_3(axpy_dp_io_out_s_3),
    .io_out_s_4(axpy_dp_io_out_s_4),
    .io_out_s_5(axpy_dp_io_out_s_5),
    .io_out_s_6(axpy_dp_io_out_s_6),
    .io_out_s_7(axpy_dp_io_out_s_7),
    .io_out_s_8(axpy_dp_io_out_s_8),
    .io_out_s_9(axpy_dp_io_out_s_9),
    .io_out_s_10(axpy_dp_io_out_s_10),
    .io_out_s_11(axpy_dp_io_out_s_11),
    .io_out_s_12(axpy_dp_io_out_s_12),
    .io_out_s_13(axpy_dp_io_out_s_13),
    .io_out_s_14(axpy_dp_io_out_s_14),
    .io_out_s_15(axpy_dp_io_out_s_15),
    .io_out_s_16(axpy_dp_io_out_s_16),
    .io_out_s_17(axpy_dp_io_out_s_17),
    .io_out_s_18(axpy_dp_io_out_s_18),
    .io_out_s_19(axpy_dp_io_out_s_19),
    .io_out_s_20(axpy_dp_io_out_s_20),
    .io_out_s_21(axpy_dp_io_out_s_21),
    .io_out_s_22(axpy_dp_io_out_s_22),
    .io_out_s_23(axpy_dp_io_out_s_23),
    .io_out_s_24(axpy_dp_io_out_s_24),
    .io_out_s_25(axpy_dp_io_out_s_25),
    .io_out_s_26(axpy_dp_io_out_s_26),
    .io_out_s_27(axpy_dp_io_out_s_27),
    .io_out_s_28(axpy_dp_io_out_s_28),
    .io_out_s_29(axpy_dp_io_out_s_29),
    .io_out_s_30(axpy_dp_io_out_s_30),
    .io_out_s_31(axpy_dp_io_out_s_31),
    .io_out_s_32(axpy_dp_io_out_s_32),
    .io_out_s_33(axpy_dp_io_out_s_33),
    .io_out_s_34(axpy_dp_io_out_s_34),
    .io_out_s_35(axpy_dp_io_out_s_35),
    .io_out_s_36(axpy_dp_io_out_s_36),
    .io_out_s_37(axpy_dp_io_out_s_37),
    .io_out_s_38(axpy_dp_io_out_s_38),
    .io_out_s_39(axpy_dp_io_out_s_39),
    .io_out_s_40(axpy_dp_io_out_s_40),
    .io_out_s_41(axpy_dp_io_out_s_41),
    .io_out_s_42(axpy_dp_io_out_s_42),
    .io_out_s_43(axpy_dp_io_out_s_43),
    .io_out_s_44(axpy_dp_io_out_s_44),
    .io_out_s_45(axpy_dp_io_out_s_45),
    .io_out_s_46(axpy_dp_io_out_s_46),
    .io_out_s_47(axpy_dp_io_out_s_47),
    .io_out_s_48(axpy_dp_io_out_s_48),
    .io_out_s_49(axpy_dp_io_out_s_49),
    .io_out_s_50(axpy_dp_io_out_s_50),
    .io_out_s_51(axpy_dp_io_out_s_51),
    .io_out_s_52(axpy_dp_io_out_s_52),
    .io_out_s_53(axpy_dp_io_out_s_53),
    .io_out_s_54(axpy_dp_io_out_s_54),
    .io_out_s_55(axpy_dp_io_out_s_55),
    .io_out_s_56(axpy_dp_io_out_s_56),
    .io_out_s_57(axpy_dp_io_out_s_57),
    .io_out_s_58(axpy_dp_io_out_s_58),
    .io_out_s_59(axpy_dp_io_out_s_59),
    .io_out_s_60(axpy_dp_io_out_s_60),
    .io_out_s_61(axpy_dp_io_out_s_61),
    .io_out_s_62(axpy_dp_io_out_s_62),
    .io_out_s_63(axpy_dp_io_out_s_63)
  );
  assign io_hh_dout = {io_hh_dout_hi,io_hh_dout_lo}; // @[hh_datapath_chisel.scala 290:28]
  assign FP_DDOT_dp_clock = io_clk;
  assign FP_DDOT_dp_reset = io_rst;
  assign FP_DDOT_dp_io_in_a_0 = ddot_din_a_reg[2047:2016]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_1 = ddot_din_a_reg[2015:1984]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_2 = ddot_din_a_reg[1983:1952]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_3 = ddot_din_a_reg[1951:1920]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_4 = ddot_din_a_reg[1919:1888]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_5 = ddot_din_a_reg[1887:1856]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_6 = ddot_din_a_reg[1855:1824]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_7 = ddot_din_a_reg[1823:1792]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_8 = ddot_din_a_reg[1791:1760]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_9 = ddot_din_a_reg[1759:1728]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_10 = ddot_din_a_reg[1727:1696]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_11 = ddot_din_a_reg[1695:1664]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_12 = ddot_din_a_reg[1663:1632]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_13 = ddot_din_a_reg[1631:1600]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_14 = ddot_din_a_reg[1599:1568]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_15 = ddot_din_a_reg[1567:1536]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_16 = ddot_din_a_reg[1535:1504]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_17 = ddot_din_a_reg[1503:1472]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_18 = ddot_din_a_reg[1471:1440]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_19 = ddot_din_a_reg[1439:1408]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_20 = ddot_din_a_reg[1407:1376]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_21 = ddot_din_a_reg[1375:1344]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_22 = ddot_din_a_reg[1343:1312]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_23 = ddot_din_a_reg[1311:1280]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_24 = ddot_din_a_reg[1279:1248]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_25 = ddot_din_a_reg[1247:1216]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_26 = ddot_din_a_reg[1215:1184]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_27 = ddot_din_a_reg[1183:1152]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_28 = ddot_din_a_reg[1151:1120]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_29 = ddot_din_a_reg[1119:1088]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_30 = ddot_din_a_reg[1087:1056]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_31 = ddot_din_a_reg[1055:1024]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_32 = ddot_din_a_reg[1023:992]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_33 = ddot_din_a_reg[991:960]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_34 = ddot_din_a_reg[959:928]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_35 = ddot_din_a_reg[927:896]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_36 = ddot_din_a_reg[895:864]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_37 = ddot_din_a_reg[863:832]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_38 = ddot_din_a_reg[831:800]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_39 = ddot_din_a_reg[799:768]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_40 = ddot_din_a_reg[767:736]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_41 = ddot_din_a_reg[735:704]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_42 = ddot_din_a_reg[703:672]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_43 = ddot_din_a_reg[671:640]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_44 = ddot_din_a_reg[639:608]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_45 = ddot_din_a_reg[607:576]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_46 = ddot_din_a_reg[575:544]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_47 = ddot_din_a_reg[543:512]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_48 = ddot_din_a_reg[511:480]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_49 = ddot_din_a_reg[479:448]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_50 = ddot_din_a_reg[447:416]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_51 = ddot_din_a_reg[415:384]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_52 = ddot_din_a_reg[383:352]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_53 = ddot_din_a_reg[351:320]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_54 = ddot_din_a_reg[319:288]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_55 = ddot_din_a_reg[287:256]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_56 = ddot_din_a_reg[255:224]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_57 = ddot_din_a_reg[223:192]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_58 = ddot_din_a_reg[191:160]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_59 = ddot_din_a_reg[159:128]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_60 = ddot_din_a_reg[127:96]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_61 = ddot_din_a_reg[95:64]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_62 = ddot_din_a_reg[63:32]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_a_63 = ddot_din_a_reg[31:0]; // @[hh_datapath_chisel.scala 251:37]
  assign FP_DDOT_dp_io_in_b_0 = ddot_din_b_reg[2047:2016]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_1 = ddot_din_b_reg[2015:1984]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_2 = ddot_din_b_reg[1983:1952]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_3 = ddot_din_b_reg[1951:1920]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_4 = ddot_din_b_reg[1919:1888]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_5 = ddot_din_b_reg[1887:1856]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_6 = ddot_din_b_reg[1855:1824]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_7 = ddot_din_b_reg[1823:1792]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_8 = ddot_din_b_reg[1791:1760]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_9 = ddot_din_b_reg[1759:1728]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_10 = ddot_din_b_reg[1727:1696]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_11 = ddot_din_b_reg[1695:1664]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_12 = ddot_din_b_reg[1663:1632]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_13 = ddot_din_b_reg[1631:1600]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_14 = ddot_din_b_reg[1599:1568]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_15 = ddot_din_b_reg[1567:1536]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_16 = ddot_din_b_reg[1535:1504]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_17 = ddot_din_b_reg[1503:1472]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_18 = ddot_din_b_reg[1471:1440]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_19 = ddot_din_b_reg[1439:1408]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_20 = ddot_din_b_reg[1407:1376]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_21 = ddot_din_b_reg[1375:1344]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_22 = ddot_din_b_reg[1343:1312]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_23 = ddot_din_b_reg[1311:1280]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_24 = ddot_din_b_reg[1279:1248]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_25 = ddot_din_b_reg[1247:1216]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_26 = ddot_din_b_reg[1215:1184]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_27 = ddot_din_b_reg[1183:1152]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_28 = ddot_din_b_reg[1151:1120]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_29 = ddot_din_b_reg[1119:1088]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_30 = ddot_din_b_reg[1087:1056]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_31 = ddot_din_b_reg[1055:1024]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_32 = ddot_din_b_reg[1023:992]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_33 = ddot_din_b_reg[991:960]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_34 = ddot_din_b_reg[959:928]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_35 = ddot_din_b_reg[927:896]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_36 = ddot_din_b_reg[895:864]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_37 = ddot_din_b_reg[863:832]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_38 = ddot_din_b_reg[831:800]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_39 = ddot_din_b_reg[799:768]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_40 = ddot_din_b_reg[767:736]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_41 = ddot_din_b_reg[735:704]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_42 = ddot_din_b_reg[703:672]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_43 = ddot_din_b_reg[671:640]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_44 = ddot_din_b_reg[639:608]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_45 = ddot_din_b_reg[607:576]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_46 = ddot_din_b_reg[575:544]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_47 = ddot_din_b_reg[543:512]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_48 = ddot_din_b_reg[511:480]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_49 = ddot_din_b_reg[479:448]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_50 = ddot_din_b_reg[447:416]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_51 = ddot_din_b_reg[415:384]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_52 = ddot_din_b_reg[383:352]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_53 = ddot_din_b_reg[351:320]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_54 = ddot_din_b_reg[319:288]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_55 = ddot_din_b_reg[287:256]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_56 = ddot_din_b_reg[255:224]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_57 = ddot_din_b_reg[223:192]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_58 = ddot_din_b_reg[191:160]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_59 = ddot_din_b_reg[159:128]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_60 = ddot_din_b_reg[127:96]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_61 = ddot_din_b_reg[95:64]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_62 = ddot_din_b_reg[63:32]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_DDOT_dp_io_in_b_63 = ddot_din_b_reg[31:0]; // @[hh_datapath_chisel.scala 252:37]
  assign FP_square_root_newfpu_clock = io_clk;
  assign FP_square_root_newfpu_reset = io_rst;
  assign FP_square_root_newfpu_io_in_a = io_d1_vld ? ddot_dout : d1_reg; // @[hh_datapath_chisel.scala 171:20 172:10 174:10]
  assign hqr5_clock = io_clk;
  assign hqr5_reset = io_rst;
  assign hqr5_io_in_a = io_d1_rdy ? x1_update : x1_reg; // @[hh_datapath_chisel.scala 183:20 184:10 186:10]
  assign hqr5_io_in_b = io_d2_vld ? d2_update : d2_reg; // @[hh_datapath_chisel.scala 189:20 190:10 192:10]
  assign hqr7_clock = io_clk;
  assign hqr7_reset = io_rst;
  assign hqr7_io_in_a = io_d3_vld ? ddot_dout : d3_reg; // @[hh_datapath_chisel.scala 177:20 178:10 180:10]
  assign FP_multiplier_10ccs_clock = io_clk;
  assign FP_multiplier_10ccs_reset = io_rst;
  assign FP_multiplier_10ccs_io_in_a = io_d5_rdy ? d4_update : d4_reg; // @[hh_datapath_chisel.scala 207:20 208:10 210:10]
  assign FP_multiplier_10ccs_io_in_b = io_tk_vld ? tk_update : tk_reg; // @[hh_datapath_chisel.scala 201:20 202:10 204:10]
  assign axpy_dp_clock = io_clk;
  assign axpy_dp_reset = io_rst;
  assign axpy_dp_io_in_a = io_d5_vld ? d5_update : d5_reg; // @[hh_datapath_chisel.scala 213:20 214:10 216:10]
  assign axpy_dp_io_in_b_0 = vk[2047:2016]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_1 = vk[2015:1984]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_2 = vk[1983:1952]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_3 = vk[1951:1920]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_4 = vk[1919:1888]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_5 = vk[1887:1856]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_6 = vk[1855:1824]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_7 = vk[1823:1792]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_8 = vk[1791:1760]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_9 = vk[1759:1728]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_10 = vk[1727:1696]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_11 = vk[1695:1664]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_12 = vk[1663:1632]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_13 = vk[1631:1600]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_14 = vk[1599:1568]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_15 = vk[1567:1536]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_16 = vk[1535:1504]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_17 = vk[1503:1472]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_18 = vk[1471:1440]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_19 = vk[1439:1408]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_20 = vk[1407:1376]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_21 = vk[1375:1344]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_22 = vk[1343:1312]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_23 = vk[1311:1280]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_24 = vk[1279:1248]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_25 = vk[1247:1216]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_26 = vk[1215:1184]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_27 = vk[1183:1152]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_28 = vk[1151:1120]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_29 = vk[1119:1088]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_30 = vk[1087:1056]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_31 = vk[1055:1024]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_32 = vk[1023:992]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_33 = vk[991:960]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_34 = vk[959:928]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_35 = vk[927:896]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_36 = vk[895:864]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_37 = vk[863:832]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_38 = vk[831:800]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_39 = vk[799:768]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_40 = vk[767:736]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_41 = vk[735:704]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_42 = vk[703:672]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_43 = vk[671:640]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_44 = vk[639:608]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_45 = vk[607:576]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_46 = vk[575:544]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_47 = vk[543:512]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_48 = vk[511:480]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_49 = vk[479:448]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_50 = vk[447:416]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_51 = vk[415:384]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_52 = vk[383:352]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_53 = vk[351:320]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_54 = vk[319:288]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_55 = vk[287:256]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_56 = vk[255:224]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_57 = vk[223:192]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_58 = vk[191:160]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_59 = vk[159:128]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_60 = vk[127:96]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_61 = vk[95:64]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_62 = vk[63:32]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_b_63 = vk[31:0]; // @[hh_datapath_chisel.scala 279:25]
  assign axpy_dp_io_in_c_0 = yj0[2047:2016]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_1 = yj0[2015:1984]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_2 = yj0[1983:1952]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_3 = yj0[1951:1920]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_4 = yj0[1919:1888]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_5 = yj0[1887:1856]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_6 = yj0[1855:1824]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_7 = yj0[1823:1792]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_8 = yj0[1791:1760]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_9 = yj0[1759:1728]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_10 = yj0[1727:1696]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_11 = yj0[1695:1664]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_12 = yj0[1663:1632]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_13 = yj0[1631:1600]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_14 = yj0[1599:1568]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_15 = yj0[1567:1536]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_16 = yj0[1535:1504]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_17 = yj0[1503:1472]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_18 = yj0[1471:1440]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_19 = yj0[1439:1408]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_20 = yj0[1407:1376]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_21 = yj0[1375:1344]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_22 = yj0[1343:1312]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_23 = yj0[1311:1280]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_24 = yj0[1279:1248]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_25 = yj0[1247:1216]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_26 = yj0[1215:1184]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_27 = yj0[1183:1152]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_28 = yj0[1151:1120]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_29 = yj0[1119:1088]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_30 = yj0[1087:1056]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_31 = yj0[1055:1024]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_32 = yj0[1023:992]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_33 = yj0[991:960]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_34 = yj0[959:928]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_35 = yj0[927:896]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_36 = yj0[895:864]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_37 = yj0[863:832]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_38 = yj0[831:800]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_39 = yj0[799:768]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_40 = yj0[767:736]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_41 = yj0[735:704]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_42 = yj0[703:672]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_43 = yj0[671:640]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_44 = yj0[639:608]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_45 = yj0[607:576]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_46 = yj0[575:544]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_47 = yj0[543:512]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_48 = yj0[511:480]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_49 = yj0[479:448]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_50 = yj0[447:416]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_51 = yj0[415:384]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_52 = yj0[383:352]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_53 = yj0[351:320]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_54 = yj0[319:288]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_55 = yj0[287:256]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_56 = yj0[255:224]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_57 = yj0[223:192]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_58 = yj0[191:160]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_59 = yj0[159:128]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_60 = yj0[127:96]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_61 = yj0[95:64]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_62 = yj0[63:32]; // @[hh_datapath_chisel.scala 280:26]
  assign axpy_dp_io_in_c_63 = yj0[31:0]; // @[hh_datapath_chisel.scala 280:26]
  always @(posedge io_clk) begin
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj0 <= 2048'h0; // @[hh_datapath_chisel.scala 64:11]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj0 <= yj_reg_4[2047:0]; // @[hh_datapath_chisel.scala 70:11]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_1 <= 116224'h0; // @[hh_datapath_chisel.scala 60:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_1 <= _yj_reg_1_T[118271:2048]; // @[hh_datapath_chisel.scala 69:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_2 <= 116224'h0; // @[hh_datapath_chisel.scala 61:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_2 <= _yj_reg_2_T_1[118271:2048]; // @[hh_datapath_chisel.scala 68:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_3 <= 116224'h0; // @[hh_datapath_chisel.scala 62:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_3 <= _yj_reg_3_T_1[118271:2048]; // @[hh_datapath_chisel.scala 67:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 59:17]
      yj_reg_4 <= 116224'h0; // @[hh_datapath_chisel.scala 63:16]
    end else if (io_yj_sft) begin // @[hh_datapath_chisel.scala 65:26]
      yj_reg_4 <= _yj_reg_4_T_1[118271:2048]; // @[hh_datapath_chisel.scala 66:16]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      ddot_din_a_reg <= 2048'h0; // @[hh_datapath_chisel.scala 110:22]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 135:20]
      ddot_din_a_reg <= io_hh_din; // @[hh_datapath_chisel.scala 136:18]
    end else if (io_d3_rdy) begin // @[hh_datapath_chisel.scala 137:26]
      if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 155:21]
        ddot_din_a_reg <= vk_update; // @[hh_datapath_chisel.scala 156:10]
      end else begin
        ddot_din_a_reg <= vk_reg; // @[hh_datapath_chisel.scala 158:10]
      end
    end else if (io_d4_rdy) begin // @[hh_datapath_chisel.scala 139:26]
      ddot_din_a_reg <= io_hh_din; // @[hh_datapath_chisel.scala 140:18]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      ddot_din_b_reg <= 2048'h0; // @[hh_datapath_chisel.scala 111:22]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 145:20]
      ddot_din_b_reg <= io_hh_din; // @[hh_datapath_chisel.scala 146:18]
    end else if (io_d3_rdy) begin // @[hh_datapath_chisel.scala 147:26]
      ddot_din_b_reg <= vk; // @[hh_datapath_chisel.scala 148:18]
    end else if (io_d4_rdy) begin // @[hh_datapath_chisel.scala 149:26]
      ddot_din_b_reg <= vk; // @[hh_datapath_chisel.scala 150:18]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      vk_reg <= 2048'h0; // @[hh_datapath_chisel.scala 112:14]
    end else if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 155:21]
      vk_reg <= vk_update; // @[hh_datapath_chisel.scala 156:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d1_reg <= 32'h0; // @[hh_datapath_chisel.scala 113:14]
    end else if (io_d1_vld) begin // @[hh_datapath_chisel.scala 171:20]
      d1_reg <= ddot_dout; // @[hh_datapath_chisel.scala 172:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d3_reg <= 32'h0; // @[hh_datapath_chisel.scala 114:14]
    end else if (io_d3_vld) begin // @[hh_datapath_chisel.scala 177:20]
      d3_reg <= ddot_dout; // @[hh_datapath_chisel.scala 178:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 162:17]
      d4_update <= 32'h0; // @[hh_datapath_chisel.scala 163:17]
    end else if (io_d4_sft) begin // @[hh_datapath_chisel.scala 165:26]
      d4_update <= d4_update_reg[31:0]; // @[hh_datapath_chisel.scala 168:17]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 115:14]
    end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 183:20]
      if (io_rst) begin // @[hh_datapath_chisel.scala 223:17]
        x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 224:17]
      end else if (io_d1_rdy) begin // @[hh_datapath_chisel.scala 225:26]
        x1_reg <= _GEN_103; // @[hh_datapath_chisel.scala 226:17]
      end else begin
        x1_reg <= 32'h0; // @[hh_datapath_chisel.scala 228:17]
      end
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d2_reg <= 32'h0; // @[hh_datapath_chisel.scala 116:14]
    end else if (io_d2_vld) begin // @[hh_datapath_chisel.scala 189:20]
      d2_reg <= d2_update; // @[hh_datapath_chisel.scala 190:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      vk1_reg <= 32'h0; // @[hh_datapath_chisel.scala 117:15]
    end else if (io_vk1_vld) begin // @[hh_datapath_chisel.scala 195:21]
      vk1_reg <= vk1_update; // @[hh_datapath_chisel.scala 196:11]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      tk_reg <= 32'h0; // @[hh_datapath_chisel.scala 118:14]
    end else if (io_tk_vld) begin // @[hh_datapath_chisel.scala 201:20]
      tk_reg <= tk_update; // @[hh_datapath_chisel.scala 202:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d4_reg <= 32'h0; // @[hh_datapath_chisel.scala 119:14]
    end else if (io_d5_rdy) begin // @[hh_datapath_chisel.scala 207:20]
      d4_reg <= d4_update; // @[hh_datapath_chisel.scala 208:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 109:18]
      d5_reg <= 32'h0; // @[hh_datapath_chisel.scala 120:14]
    end else if (io_d5_vld) begin // @[hh_datapath_chisel.scala 213:20]
      d5_reg <= d5_update; // @[hh_datapath_chisel.scala 214:10]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 162:17]
      d4_update_reg <= 4064'h0; // @[hh_datapath_chisel.scala 164:21]
    end else if (io_d4_sft) begin // @[hh_datapath_chisel.scala 165:26]
      d4_update_reg <= _d4_update_reg_T[4095:32]; // @[hh_datapath_chisel.scala 167:21]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_0 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_0 <= axpy_dp_io_out_s_63; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_1 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_1 <= axpy_dp_io_out_s_62; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_2 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_2 <= axpy_dp_io_out_s_61; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_3 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_3 <= axpy_dp_io_out_s_60; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_4 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_4 <= axpy_dp_io_out_s_59; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_5 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_5 <= axpy_dp_io_out_s_58; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_6 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_6 <= axpy_dp_io_out_s_57; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_7 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_7 <= axpy_dp_io_out_s_56; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_8 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_8 <= axpy_dp_io_out_s_55; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_9 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_9 <= axpy_dp_io_out_s_54; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_10 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_10 <= axpy_dp_io_out_s_53; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_11 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_11 <= axpy_dp_io_out_s_52; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_12 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_12 <= axpy_dp_io_out_s_51; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_13 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_13 <= axpy_dp_io_out_s_50; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_14 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_14 <= axpy_dp_io_out_s_49; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_15 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_15 <= axpy_dp_io_out_s_48; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_16 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_16 <= axpy_dp_io_out_s_47; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_17 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_17 <= axpy_dp_io_out_s_46; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_18 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_18 <= axpy_dp_io_out_s_45; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_19 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_19 <= axpy_dp_io_out_s_44; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_20 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_20 <= axpy_dp_io_out_s_43; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_21 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_21 <= axpy_dp_io_out_s_42; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_22 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_22 <= axpy_dp_io_out_s_41; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_23 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_23 <= axpy_dp_io_out_s_40; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_24 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_24 <= axpy_dp_io_out_s_39; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_25 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_25 <= axpy_dp_io_out_s_38; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_26 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_26 <= axpy_dp_io_out_s_37; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_27 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_27 <= axpy_dp_io_out_s_36; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_28 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_28 <= axpy_dp_io_out_s_35; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_29 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_29 <= axpy_dp_io_out_s_34; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_30 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_30 <= axpy_dp_io_out_s_33; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_31 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_31 <= axpy_dp_io_out_s_32; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_32 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_32 <= axpy_dp_io_out_s_31; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_33 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_33 <= axpy_dp_io_out_s_30; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_34 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_34 <= axpy_dp_io_out_s_29; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_35 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_35 <= axpy_dp_io_out_s_28; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_36 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_36 <= axpy_dp_io_out_s_27; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_37 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_37 <= axpy_dp_io_out_s_26; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_38 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_38 <= axpy_dp_io_out_s_25; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_39 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_39 <= axpy_dp_io_out_s_24; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_40 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_40 <= axpy_dp_io_out_s_23; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_41 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_41 <= axpy_dp_io_out_s_22; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_42 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_42 <= axpy_dp_io_out_s_21; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_43 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_43 <= axpy_dp_io_out_s_20; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_44 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_44 <= axpy_dp_io_out_s_19; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_45 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_45 <= axpy_dp_io_out_s_18; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_46 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_46 <= axpy_dp_io_out_s_17; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_47 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_47 <= axpy_dp_io_out_s_16; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_48 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_48 <= axpy_dp_io_out_s_15; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_49 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_49 <= axpy_dp_io_out_s_14; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_50 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_50 <= axpy_dp_io_out_s_13; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_51 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_51 <= axpy_dp_io_out_s_12; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_52 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_52 <= axpy_dp_io_out_s_11; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_53 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_53 <= axpy_dp_io_out_s_10; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_54 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_54 <= axpy_dp_io_out_s_9; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_55 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_55 <= axpy_dp_io_out_s_8; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_56 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_56 <= axpy_dp_io_out_s_7; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_57 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_57 <= axpy_dp_io_out_s_6; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_58 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_58 <= axpy_dp_io_out_s_5; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_59 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_59 <= axpy_dp_io_out_s_4; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_60 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_60 <= axpy_dp_io_out_s_3; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_61 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_61 <= axpy_dp_io_out_s_2; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_62 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_62 <= axpy_dp_io_out_s_1; // @[hh_datapath_chisel.scala 288:36]
    end
    if (io_rst) begin // @[hh_datapath_chisel.scala 283:16]
      myAxpyVec_63 <= 32'h0; // @[hh_datapath_chisel.scala 285:36]
    end else begin
      myAxpyVec_63 <= axpy_dp_io_out_s_0; // @[hh_datapath_chisel.scala 288:36]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {64{`RANDOM}};
  yj0 = _RAND_0[2047:0];
  _RAND_1 = {3632{`RANDOM}};
  yj_reg_1 = _RAND_1[116223:0];
  _RAND_2 = {3632{`RANDOM}};
  yj_reg_2 = _RAND_2[116223:0];
  _RAND_3 = {3632{`RANDOM}};
  yj_reg_3 = _RAND_3[116223:0];
  _RAND_4 = {3632{`RANDOM}};
  yj_reg_4 = _RAND_4[116223:0];
  _RAND_5 = {64{`RANDOM}};
  ddot_din_a_reg = _RAND_5[2047:0];
  _RAND_6 = {64{`RANDOM}};
  ddot_din_b_reg = _RAND_6[2047:0];
  _RAND_7 = {64{`RANDOM}};
  vk_reg = _RAND_7[2047:0];
  _RAND_8 = {1{`RANDOM}};
  d1_reg = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  d3_reg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  d4_update = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  x1_reg = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  d2_reg = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  vk1_reg = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  tk_reg = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  d4_reg = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  d5_reg = _RAND_16[31:0];
  _RAND_17 = {127{`RANDOM}};
  d4_update_reg = _RAND_17[4063:0];
  _RAND_18 = {1{`RANDOM}};
  myAxpyVec_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  myAxpyVec_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  myAxpyVec_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  myAxpyVec_3 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  myAxpyVec_4 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  myAxpyVec_5 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  myAxpyVec_6 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  myAxpyVec_7 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  myAxpyVec_8 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  myAxpyVec_9 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  myAxpyVec_10 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  myAxpyVec_11 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  myAxpyVec_12 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  myAxpyVec_13 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  myAxpyVec_14 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  myAxpyVec_15 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  myAxpyVec_16 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  myAxpyVec_17 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  myAxpyVec_18 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  myAxpyVec_19 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  myAxpyVec_20 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  myAxpyVec_21 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  myAxpyVec_22 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  myAxpyVec_23 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  myAxpyVec_24 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  myAxpyVec_25 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  myAxpyVec_26 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  myAxpyVec_27 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  myAxpyVec_28 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  myAxpyVec_29 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  myAxpyVec_30 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  myAxpyVec_31 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  myAxpyVec_32 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  myAxpyVec_33 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  myAxpyVec_34 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  myAxpyVec_35 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  myAxpyVec_36 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  myAxpyVec_37 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  myAxpyVec_38 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  myAxpyVec_39 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  myAxpyVec_40 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  myAxpyVec_41 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  myAxpyVec_42 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  myAxpyVec_43 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  myAxpyVec_44 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  myAxpyVec_45 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  myAxpyVec_46 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  myAxpyVec_47 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  myAxpyVec_48 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  myAxpyVec_49 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  myAxpyVec_50 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  myAxpyVec_51 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  myAxpyVec_52 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  myAxpyVec_53 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  myAxpyVec_54 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  myAxpyVec_55 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  myAxpyVec_56 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  myAxpyVec_57 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  myAxpyVec_58 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  myAxpyVec_59 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  myAxpyVec_60 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  myAxpyVec_61 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  myAxpyVec_62 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  myAxpyVec_63 = _RAND_81[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module hh_core(
  input           io_clk,
  input           io_rst,
  input  [15:0]   io_hh_cnt,
  input           io_d1_rdy,
  input           io_d1_vld,
  input           io_d2_vld,
  input           io_vk1_vld,
  input           io_d3_rdy,
  input           io_d3_vld,
  input           io_tk_vld,
  input           io_d4_rdy,
  input           io_d5_rdy,
  input           io_d5_vld,
  input           io_yj_sft,
  input           io_d4_sft,
  input           io_hh_st,
  input           io_dmx0_mem_ena,
  input  [127:0]  io_dmx0_mem_wea,
  input  [4:0]    io_dmx0_mem_addra,
  input  [1023:0] io_dmx0_mem_dina,
  input           io_dmx0_mem_enb,
  input  [4:0]    io_dmx0_mem_addrb,
  output [1023:0] io_dmx0_mem_doutb,
  input           io_dmx1_mem_ena,
  input  [127:0]  io_dmx1_mem_wea,
  input  [4:0]    io_dmx1_mem_addra,
  input  [1023:0] io_dmx1_mem_dina,
  input           io_dmx1_mem_enb,
  input  [4:0]    io_dmx1_mem_addrb,
  output [1023:0] io_dmx1_mem_doutb,
  input           io_rtri_mem_ena,
  input  [127:0]  io_rtri_mem_wea,
  input  [4:0]    io_rtri_mem_addra,
  input  [1023:0] io_rtri_mem_dina,
  input           io_rtri_mem_enb,
  input  [4:0]    io_rtri_mem_addrb,
  output [1023:0] io_rtri_mem_doutb,
  output [2047:0] io_hh_dout
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [2047:0] _RAND_2;
  reg [2047:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  simple_dual_io_clka; // @[hh_core.scala 163:31]
  wire  simple_dual_io_clkb; // @[hh_core.scala 163:31]
  wire  simple_dual_io_ena; // @[hh_core.scala 163:31]
  wire  simple_dual_io_enb; // @[hh_core.scala 163:31]
  wire [127:0] simple_dual_io_wea; // @[hh_core.scala 163:31]
  wire [4:0] simple_dual_io_addra; // @[hh_core.scala 163:31]
  wire [4:0] simple_dual_io_addrb; // @[hh_core.scala 163:31]
  wire [1023:0] simple_dual_io_dina; // @[hh_core.scala 163:31]
  wire [1023:0] simple_dual_io_doutb; // @[hh_core.scala 163:31]
  wire  simple_dual_1_io_clka; // @[hh_core.scala 175:31]
  wire  simple_dual_1_io_clkb; // @[hh_core.scala 175:31]
  wire  simple_dual_1_io_ena; // @[hh_core.scala 175:31]
  wire  simple_dual_1_io_enb; // @[hh_core.scala 175:31]
  wire [127:0] simple_dual_1_io_wea; // @[hh_core.scala 175:31]
  wire [4:0] simple_dual_1_io_addra; // @[hh_core.scala 175:31]
  wire [4:0] simple_dual_1_io_addrb; // @[hh_core.scala 175:31]
  wire [1023:0] simple_dual_1_io_dina; // @[hh_core.scala 175:31]
  wire [1023:0] simple_dual_1_io_doutb; // @[hh_core.scala 175:31]
  wire  simple_dual_2_io_clka; // @[hh_core.scala 186:31]
  wire  simple_dual_2_io_clkb; // @[hh_core.scala 186:31]
  wire  simple_dual_2_io_ena; // @[hh_core.scala 186:31]
  wire  simple_dual_2_io_enb; // @[hh_core.scala 186:31]
  wire [127:0] simple_dual_2_io_wea; // @[hh_core.scala 186:31]
  wire [4:0] simple_dual_2_io_addra; // @[hh_core.scala 186:31]
  wire [4:0] simple_dual_2_io_addrb; // @[hh_core.scala 186:31]
  wire [1023:0] simple_dual_2_io_dina; // @[hh_core.scala 186:31]
  wire [1023:0] simple_dual_2_io_doutb; // @[hh_core.scala 186:31]
  wire  u_hh_datapath_io_clk; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_rst; // @[hh_core.scala 197:38]
  wire [15:0] u_hh_datapath_io_hh_cnt; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d1_rdy; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d1_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d2_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_vk1_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d3_rdy; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d3_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_tk_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d4_rdy; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d5_rdy; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d5_vld; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_yj_sft; // @[hh_core.scala 197:38]
  wire  u_hh_datapath_io_d4_sft; // @[hh_core.scala 197:38]
  wire [2047:0] u_hh_datapath_io_hh_din; // @[hh_core.scala 197:38]
  wire [2047:0] u_hh_datapath_io_hh_dout; // @[hh_core.scala 197:38]
  reg  hh0_din_rdy; // @[hh_core.scala 79:34]
  reg  hh1_din_rdy; // @[hh_core.scala 80:34]
  reg [2047:0] hh_din_reg; // @[hh_core.scala 82:33]
  reg [2047:0] hh_din; // @[hh_core.scala 85:29]
  wire  _T = hh0_din_rdy | hh1_din_rdy; // @[hh_core.scala 100:30]
  wire [16:0] _myTriMemVec2_31_T = {{1'd0}, io_hh_cnt}; // @[hh_core.scala 127:74]
  wire [31:0] myTriMemVec_31 = io_rtri_mem_doutb[31:0]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_30 = io_rtri_mem_doutb[63:32]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_29 = io_rtri_mem_doutb[95:64]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_28 = io_rtri_mem_doutb[127:96]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_27 = io_rtri_mem_doutb[159:128]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_26 = io_rtri_mem_doutb[191:160]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_25 = io_rtri_mem_doutb[223:192]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_24 = io_rtri_mem_doutb[255:224]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_23 = io_rtri_mem_doutb[287:256]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_22 = io_rtri_mem_doutb[319:288]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_21 = io_rtri_mem_doutb[351:320]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_20 = io_rtri_mem_doutb[383:352]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_19 = io_rtri_mem_doutb[415:384]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_18 = io_rtri_mem_doutb[447:416]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_17 = io_rtri_mem_doutb[479:448]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_16 = io_rtri_mem_doutb[511:480]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_15 = io_rtri_mem_doutb[543:512]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_14 = io_rtri_mem_doutb[575:544]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_13 = io_rtri_mem_doutb[607:576]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_12 = io_rtri_mem_doutb[639:608]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_11 = io_rtri_mem_doutb[671:640]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_10 = io_rtri_mem_doutb[703:672]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_9 = io_rtri_mem_doutb[735:704]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_8 = io_rtri_mem_doutb[767:736]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_7 = io_rtri_mem_doutb[799:768]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_6 = io_rtri_mem_doutb[831:800]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_5 = io_rtri_mem_doutb[863:832]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_4 = io_rtri_mem_doutb[895:864]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_3 = io_rtri_mem_doutb[927:896]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_2 = io_rtri_mem_doutb[959:928]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_1 = io_rtri_mem_doutb[991:960]; // @[hh_core.scala 122:52]
  wire [31:0] myTriMemVec_0 = io_rtri_mem_doutb[1023:992]; // @[hh_core.scala 122:52]
  wire [31:0] _GEN_8 = 5'h1 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_9 = 5'h2 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_2 : _GEN_8; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_10 = 5'h3 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_3 : _GEN_9; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_11 = 5'h4 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_4 : _GEN_10; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_12 = 5'h5 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_5 : _GEN_11; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_13 = 5'h6 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_6 : _GEN_12; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_14 = 5'h7 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_7 : _GEN_13; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_15 = 5'h8 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_8 : _GEN_14; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_16 = 5'h9 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_9 : _GEN_15; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_17 = 5'ha == _myTriMemVec2_31_T[4:0] ? myTriMemVec_10 : _GEN_16; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_18 = 5'hb == _myTriMemVec2_31_T[4:0] ? myTriMemVec_11 : _GEN_17; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_19 = 5'hc == _myTriMemVec2_31_T[4:0] ? myTriMemVec_12 : _GEN_18; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_20 = 5'hd == _myTriMemVec2_31_T[4:0] ? myTriMemVec_13 : _GEN_19; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_21 = 5'he == _myTriMemVec2_31_T[4:0] ? myTriMemVec_14 : _GEN_20; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_22 = 5'hf == _myTriMemVec2_31_T[4:0] ? myTriMemVec_15 : _GEN_21; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_23 = 5'h10 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_16 : _GEN_22; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_24 = 5'h11 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_17 : _GEN_23; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_25 = 5'h12 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_18 : _GEN_24; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_26 = 5'h13 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_19 : _GEN_25; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_27 = 5'h14 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_20 : _GEN_26; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_28 = 5'h15 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_21 : _GEN_27; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_29 = 5'h16 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_22 : _GEN_28; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_30 = 5'h17 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_23 : _GEN_29; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_31 = 5'h18 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_24 : _GEN_30; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_32 = 5'h19 == _myTriMemVec2_31_T[4:0] ? myTriMemVec_25 : _GEN_31; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_33 = 5'h1a == _myTriMemVec2_31_T[4:0] ? myTriMemVec_26 : _GEN_32; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_34 = 5'h1b == _myTriMemVec2_31_T[4:0] ? myTriMemVec_27 : _GEN_33; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_35 = 5'h1c == _myTriMemVec2_31_T[4:0] ? myTriMemVec_28 : _GEN_34; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_36 = 5'h1d == _myTriMemVec2_31_T[4:0] ? myTriMemVec_29 : _GEN_35; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_37 = 5'h1e == _myTriMemVec2_31_T[4:0] ? myTriMemVec_30 : _GEN_36; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_31 = 5'h1f == _myTriMemVec2_31_T[4:0] ? myTriMemVec_31 : _GEN_37; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_30_T_1 = 16'h1 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_40 = 5'h1 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_41 = 5'h2 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_2 : _GEN_40; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_42 = 5'h3 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_3 : _GEN_41; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_43 = 5'h4 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_4 : _GEN_42; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_44 = 5'h5 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_5 : _GEN_43; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_45 = 5'h6 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_6 : _GEN_44; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_46 = 5'h7 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_7 : _GEN_45; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_47 = 5'h8 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_8 : _GEN_46; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_48 = 5'h9 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_9 : _GEN_47; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_49 = 5'ha == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_10 : _GEN_48; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_50 = 5'hb == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_11 : _GEN_49; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_51 = 5'hc == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_12 : _GEN_50; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_52 = 5'hd == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_13 : _GEN_51; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_53 = 5'he == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_14 : _GEN_52; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_54 = 5'hf == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_15 : _GEN_53; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_55 = 5'h10 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_16 : _GEN_54; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_56 = 5'h11 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_17 : _GEN_55; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_57 = 5'h12 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_18 : _GEN_56; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_58 = 5'h13 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_19 : _GEN_57; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_59 = 5'h14 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_20 : _GEN_58; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_60 = 5'h15 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_21 : _GEN_59; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_61 = 5'h16 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_22 : _GEN_60; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_62 = 5'h17 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_23 : _GEN_61; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_63 = 5'h18 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_24 : _GEN_62; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_64 = 5'h19 == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_25 : _GEN_63; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_65 = 5'h1a == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_26 : _GEN_64; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_66 = 5'h1b == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_27 : _GEN_65; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_67 = 5'h1c == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_28 : _GEN_66; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_68 = 5'h1d == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_29 : _GEN_67; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_69 = 5'h1e == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_30 : _GEN_68; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_30 = 5'h1f == _myTriMemVec2_30_T_1[4:0] ? myTriMemVec_31 : _GEN_69; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_29_T_1 = 16'h2 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_72 = 5'h1 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_73 = 5'h2 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_2 : _GEN_72; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_74 = 5'h3 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_3 : _GEN_73; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_75 = 5'h4 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_4 : _GEN_74; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_76 = 5'h5 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_5 : _GEN_75; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_77 = 5'h6 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_6 : _GEN_76; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_78 = 5'h7 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_7 : _GEN_77; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_79 = 5'h8 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_8 : _GEN_78; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_80 = 5'h9 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_9 : _GEN_79; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_81 = 5'ha == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_10 : _GEN_80; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_82 = 5'hb == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_11 : _GEN_81; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_83 = 5'hc == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_12 : _GEN_82; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_84 = 5'hd == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_13 : _GEN_83; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_85 = 5'he == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_14 : _GEN_84; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_86 = 5'hf == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_15 : _GEN_85; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_87 = 5'h10 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_16 : _GEN_86; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_88 = 5'h11 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_17 : _GEN_87; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_89 = 5'h12 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_18 : _GEN_88; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_90 = 5'h13 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_19 : _GEN_89; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_91 = 5'h14 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_20 : _GEN_90; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_92 = 5'h15 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_21 : _GEN_91; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_93 = 5'h16 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_22 : _GEN_92; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_94 = 5'h17 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_23 : _GEN_93; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_95 = 5'h18 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_24 : _GEN_94; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_96 = 5'h19 == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_25 : _GEN_95; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_97 = 5'h1a == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_26 : _GEN_96; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_98 = 5'h1b == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_27 : _GEN_97; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_99 = 5'h1c == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_28 : _GEN_98; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_100 = 5'h1d == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_29 : _GEN_99; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_101 = 5'h1e == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_30 : _GEN_100; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_29 = 5'h1f == _myTriMemVec2_29_T_1[4:0] ? myTriMemVec_31 : _GEN_101; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_28_T_1 = 16'h3 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_104 = 5'h1 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_105 = 5'h2 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_2 : _GEN_104; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_106 = 5'h3 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_3 : _GEN_105; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_107 = 5'h4 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_4 : _GEN_106; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_108 = 5'h5 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_5 : _GEN_107; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_109 = 5'h6 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_6 : _GEN_108; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_110 = 5'h7 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_7 : _GEN_109; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_111 = 5'h8 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_8 : _GEN_110; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_112 = 5'h9 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_9 : _GEN_111; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_113 = 5'ha == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_10 : _GEN_112; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_114 = 5'hb == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_11 : _GEN_113; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_115 = 5'hc == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_12 : _GEN_114; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_116 = 5'hd == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_13 : _GEN_115; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_117 = 5'he == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_14 : _GEN_116; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_118 = 5'hf == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_15 : _GEN_117; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_119 = 5'h10 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_16 : _GEN_118; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_120 = 5'h11 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_17 : _GEN_119; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_121 = 5'h12 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_18 : _GEN_120; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_122 = 5'h13 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_19 : _GEN_121; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_123 = 5'h14 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_20 : _GEN_122; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_124 = 5'h15 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_21 : _GEN_123; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_125 = 5'h16 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_22 : _GEN_124; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_126 = 5'h17 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_23 : _GEN_125; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_127 = 5'h18 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_24 : _GEN_126; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_128 = 5'h19 == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_25 : _GEN_127; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_129 = 5'h1a == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_26 : _GEN_128; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_130 = 5'h1b == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_27 : _GEN_129; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_131 = 5'h1c == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_28 : _GEN_130; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_132 = 5'h1d == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_29 : _GEN_131; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_133 = 5'h1e == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_30 : _GEN_132; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_28 = 5'h1f == _myTriMemVec2_28_T_1[4:0] ? myTriMemVec_31 : _GEN_133; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_27_T_1 = 16'h4 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_136 = 5'h1 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_137 = 5'h2 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_2 : _GEN_136; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_138 = 5'h3 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_3 : _GEN_137; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_139 = 5'h4 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_4 : _GEN_138; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_140 = 5'h5 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_5 : _GEN_139; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_141 = 5'h6 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_6 : _GEN_140; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_142 = 5'h7 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_7 : _GEN_141; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_143 = 5'h8 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_8 : _GEN_142; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_144 = 5'h9 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_9 : _GEN_143; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_145 = 5'ha == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_10 : _GEN_144; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_146 = 5'hb == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_11 : _GEN_145; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_147 = 5'hc == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_12 : _GEN_146; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_148 = 5'hd == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_13 : _GEN_147; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_149 = 5'he == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_14 : _GEN_148; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_150 = 5'hf == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_15 : _GEN_149; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_151 = 5'h10 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_16 : _GEN_150; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_152 = 5'h11 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_17 : _GEN_151; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_153 = 5'h12 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_18 : _GEN_152; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_154 = 5'h13 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_19 : _GEN_153; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_155 = 5'h14 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_20 : _GEN_154; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_156 = 5'h15 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_21 : _GEN_155; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_157 = 5'h16 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_22 : _GEN_156; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_158 = 5'h17 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_23 : _GEN_157; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_159 = 5'h18 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_24 : _GEN_158; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_160 = 5'h19 == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_25 : _GEN_159; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_161 = 5'h1a == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_26 : _GEN_160; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_162 = 5'h1b == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_27 : _GEN_161; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_163 = 5'h1c == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_28 : _GEN_162; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_164 = 5'h1d == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_29 : _GEN_163; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_165 = 5'h1e == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_30 : _GEN_164; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_27 = 5'h1f == _myTriMemVec2_27_T_1[4:0] ? myTriMemVec_31 : _GEN_165; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_26_T_1 = 16'h5 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_168 = 5'h1 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_169 = 5'h2 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_2 : _GEN_168; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_170 = 5'h3 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_3 : _GEN_169; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_171 = 5'h4 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_4 : _GEN_170; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_172 = 5'h5 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_5 : _GEN_171; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_173 = 5'h6 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_6 : _GEN_172; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_174 = 5'h7 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_7 : _GEN_173; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_175 = 5'h8 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_8 : _GEN_174; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_176 = 5'h9 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_9 : _GEN_175; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_177 = 5'ha == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_10 : _GEN_176; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_178 = 5'hb == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_11 : _GEN_177; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_179 = 5'hc == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_12 : _GEN_178; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_180 = 5'hd == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_13 : _GEN_179; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_181 = 5'he == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_14 : _GEN_180; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_182 = 5'hf == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_15 : _GEN_181; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_183 = 5'h10 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_16 : _GEN_182; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_184 = 5'h11 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_17 : _GEN_183; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_185 = 5'h12 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_18 : _GEN_184; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_186 = 5'h13 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_19 : _GEN_185; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_187 = 5'h14 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_20 : _GEN_186; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_188 = 5'h15 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_21 : _GEN_187; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_189 = 5'h16 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_22 : _GEN_188; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_190 = 5'h17 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_23 : _GEN_189; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_191 = 5'h18 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_24 : _GEN_190; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_192 = 5'h19 == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_25 : _GEN_191; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_193 = 5'h1a == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_26 : _GEN_192; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_194 = 5'h1b == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_27 : _GEN_193; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_195 = 5'h1c == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_28 : _GEN_194; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_196 = 5'h1d == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_29 : _GEN_195; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_197 = 5'h1e == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_30 : _GEN_196; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_26 = 5'h1f == _myTriMemVec2_26_T_1[4:0] ? myTriMemVec_31 : _GEN_197; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_25_T_1 = 16'h6 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_200 = 5'h1 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_201 = 5'h2 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_2 : _GEN_200; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_202 = 5'h3 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_3 : _GEN_201; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_203 = 5'h4 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_4 : _GEN_202; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_204 = 5'h5 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_5 : _GEN_203; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_205 = 5'h6 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_6 : _GEN_204; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_206 = 5'h7 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_7 : _GEN_205; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_207 = 5'h8 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_8 : _GEN_206; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_208 = 5'h9 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_9 : _GEN_207; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_209 = 5'ha == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_10 : _GEN_208; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_210 = 5'hb == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_11 : _GEN_209; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_211 = 5'hc == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_12 : _GEN_210; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_212 = 5'hd == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_13 : _GEN_211; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_213 = 5'he == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_14 : _GEN_212; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_214 = 5'hf == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_15 : _GEN_213; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_215 = 5'h10 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_16 : _GEN_214; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_216 = 5'h11 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_17 : _GEN_215; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_217 = 5'h12 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_18 : _GEN_216; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_218 = 5'h13 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_19 : _GEN_217; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_219 = 5'h14 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_20 : _GEN_218; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_220 = 5'h15 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_21 : _GEN_219; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_221 = 5'h16 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_22 : _GEN_220; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_222 = 5'h17 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_23 : _GEN_221; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_223 = 5'h18 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_24 : _GEN_222; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_224 = 5'h19 == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_25 : _GEN_223; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_225 = 5'h1a == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_26 : _GEN_224; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_226 = 5'h1b == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_27 : _GEN_225; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_227 = 5'h1c == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_28 : _GEN_226; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_228 = 5'h1d == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_29 : _GEN_227; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_229 = 5'h1e == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_30 : _GEN_228; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_25 = 5'h1f == _myTriMemVec2_25_T_1[4:0] ? myTriMemVec_31 : _GEN_229; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_24_T_1 = 16'h7 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_232 = 5'h1 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_233 = 5'h2 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_2 : _GEN_232; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_234 = 5'h3 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_3 : _GEN_233; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_235 = 5'h4 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_4 : _GEN_234; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_236 = 5'h5 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_5 : _GEN_235; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_237 = 5'h6 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_6 : _GEN_236; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_238 = 5'h7 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_7 : _GEN_237; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_239 = 5'h8 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_8 : _GEN_238; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_240 = 5'h9 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_9 : _GEN_239; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_241 = 5'ha == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_10 : _GEN_240; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_242 = 5'hb == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_11 : _GEN_241; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_243 = 5'hc == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_12 : _GEN_242; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_244 = 5'hd == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_13 : _GEN_243; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_245 = 5'he == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_14 : _GEN_244; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_246 = 5'hf == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_15 : _GEN_245; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_247 = 5'h10 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_16 : _GEN_246; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_248 = 5'h11 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_17 : _GEN_247; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_249 = 5'h12 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_18 : _GEN_248; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_250 = 5'h13 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_19 : _GEN_249; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_251 = 5'h14 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_20 : _GEN_250; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_252 = 5'h15 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_21 : _GEN_251; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_253 = 5'h16 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_22 : _GEN_252; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_254 = 5'h17 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_23 : _GEN_253; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_255 = 5'h18 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_24 : _GEN_254; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_256 = 5'h19 == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_25 : _GEN_255; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_257 = 5'h1a == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_26 : _GEN_256; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_258 = 5'h1b == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_27 : _GEN_257; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_259 = 5'h1c == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_28 : _GEN_258; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_260 = 5'h1d == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_29 : _GEN_259; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_261 = 5'h1e == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_30 : _GEN_260; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_24 = 5'h1f == _myTriMemVec2_24_T_1[4:0] ? myTriMemVec_31 : _GEN_261; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_23_T_1 = 16'h8 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_264 = 5'h1 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_265 = 5'h2 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_2 : _GEN_264; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_266 = 5'h3 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_3 : _GEN_265; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_267 = 5'h4 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_4 : _GEN_266; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_268 = 5'h5 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_5 : _GEN_267; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_269 = 5'h6 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_6 : _GEN_268; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_270 = 5'h7 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_7 : _GEN_269; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_271 = 5'h8 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_8 : _GEN_270; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_272 = 5'h9 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_9 : _GEN_271; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_273 = 5'ha == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_10 : _GEN_272; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_274 = 5'hb == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_11 : _GEN_273; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_275 = 5'hc == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_12 : _GEN_274; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_276 = 5'hd == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_13 : _GEN_275; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_277 = 5'he == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_14 : _GEN_276; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_278 = 5'hf == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_15 : _GEN_277; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_279 = 5'h10 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_16 : _GEN_278; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_280 = 5'h11 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_17 : _GEN_279; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_281 = 5'h12 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_18 : _GEN_280; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_282 = 5'h13 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_19 : _GEN_281; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_283 = 5'h14 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_20 : _GEN_282; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_284 = 5'h15 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_21 : _GEN_283; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_285 = 5'h16 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_22 : _GEN_284; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_286 = 5'h17 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_23 : _GEN_285; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_287 = 5'h18 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_24 : _GEN_286; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_288 = 5'h19 == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_25 : _GEN_287; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_289 = 5'h1a == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_26 : _GEN_288; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_290 = 5'h1b == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_27 : _GEN_289; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_291 = 5'h1c == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_28 : _GEN_290; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_292 = 5'h1d == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_29 : _GEN_291; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_293 = 5'h1e == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_30 : _GEN_292; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_23 = 5'h1f == _myTriMemVec2_23_T_1[4:0] ? myTriMemVec_31 : _GEN_293; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_22_T_1 = 16'h9 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_296 = 5'h1 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_297 = 5'h2 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_2 : _GEN_296; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_298 = 5'h3 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_3 : _GEN_297; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_299 = 5'h4 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_4 : _GEN_298; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_300 = 5'h5 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_5 : _GEN_299; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_301 = 5'h6 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_6 : _GEN_300; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_302 = 5'h7 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_7 : _GEN_301; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_303 = 5'h8 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_8 : _GEN_302; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_304 = 5'h9 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_9 : _GEN_303; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_305 = 5'ha == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_10 : _GEN_304; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_306 = 5'hb == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_11 : _GEN_305; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_307 = 5'hc == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_12 : _GEN_306; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_308 = 5'hd == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_13 : _GEN_307; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_309 = 5'he == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_14 : _GEN_308; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_310 = 5'hf == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_15 : _GEN_309; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_311 = 5'h10 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_16 : _GEN_310; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_312 = 5'h11 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_17 : _GEN_311; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_313 = 5'h12 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_18 : _GEN_312; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_314 = 5'h13 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_19 : _GEN_313; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_315 = 5'h14 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_20 : _GEN_314; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_316 = 5'h15 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_21 : _GEN_315; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_317 = 5'h16 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_22 : _GEN_316; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_318 = 5'h17 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_23 : _GEN_317; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_319 = 5'h18 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_24 : _GEN_318; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_320 = 5'h19 == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_25 : _GEN_319; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_321 = 5'h1a == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_26 : _GEN_320; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_322 = 5'h1b == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_27 : _GEN_321; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_323 = 5'h1c == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_28 : _GEN_322; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_324 = 5'h1d == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_29 : _GEN_323; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_325 = 5'h1e == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_30 : _GEN_324; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_22 = 5'h1f == _myTriMemVec2_22_T_1[4:0] ? myTriMemVec_31 : _GEN_325; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_21_T_1 = 16'ha + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_328 = 5'h1 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_329 = 5'h2 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_2 : _GEN_328; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_330 = 5'h3 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_3 : _GEN_329; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_331 = 5'h4 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_4 : _GEN_330; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_332 = 5'h5 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_5 : _GEN_331; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_333 = 5'h6 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_6 : _GEN_332; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_334 = 5'h7 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_7 : _GEN_333; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_335 = 5'h8 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_8 : _GEN_334; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_336 = 5'h9 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_9 : _GEN_335; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_337 = 5'ha == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_10 : _GEN_336; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_338 = 5'hb == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_11 : _GEN_337; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_339 = 5'hc == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_12 : _GEN_338; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_340 = 5'hd == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_13 : _GEN_339; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_341 = 5'he == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_14 : _GEN_340; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_342 = 5'hf == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_15 : _GEN_341; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_343 = 5'h10 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_16 : _GEN_342; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_344 = 5'h11 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_17 : _GEN_343; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_345 = 5'h12 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_18 : _GEN_344; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_346 = 5'h13 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_19 : _GEN_345; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_347 = 5'h14 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_20 : _GEN_346; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_348 = 5'h15 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_21 : _GEN_347; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_349 = 5'h16 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_22 : _GEN_348; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_350 = 5'h17 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_23 : _GEN_349; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_351 = 5'h18 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_24 : _GEN_350; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_352 = 5'h19 == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_25 : _GEN_351; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_353 = 5'h1a == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_26 : _GEN_352; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_354 = 5'h1b == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_27 : _GEN_353; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_355 = 5'h1c == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_28 : _GEN_354; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_356 = 5'h1d == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_29 : _GEN_355; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_357 = 5'h1e == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_30 : _GEN_356; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_21 = 5'h1f == _myTriMemVec2_21_T_1[4:0] ? myTriMemVec_31 : _GEN_357; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_20_T_1 = 16'hb + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_360 = 5'h1 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_361 = 5'h2 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_2 : _GEN_360; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_362 = 5'h3 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_3 : _GEN_361; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_363 = 5'h4 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_4 : _GEN_362; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_364 = 5'h5 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_5 : _GEN_363; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_365 = 5'h6 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_6 : _GEN_364; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_366 = 5'h7 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_7 : _GEN_365; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_367 = 5'h8 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_8 : _GEN_366; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_368 = 5'h9 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_9 : _GEN_367; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_369 = 5'ha == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_10 : _GEN_368; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_370 = 5'hb == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_11 : _GEN_369; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_371 = 5'hc == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_12 : _GEN_370; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_372 = 5'hd == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_13 : _GEN_371; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_373 = 5'he == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_14 : _GEN_372; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_374 = 5'hf == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_15 : _GEN_373; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_375 = 5'h10 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_16 : _GEN_374; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_376 = 5'h11 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_17 : _GEN_375; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_377 = 5'h12 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_18 : _GEN_376; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_378 = 5'h13 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_19 : _GEN_377; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_379 = 5'h14 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_20 : _GEN_378; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_380 = 5'h15 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_21 : _GEN_379; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_381 = 5'h16 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_22 : _GEN_380; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_382 = 5'h17 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_23 : _GEN_381; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_383 = 5'h18 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_24 : _GEN_382; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_384 = 5'h19 == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_25 : _GEN_383; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_385 = 5'h1a == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_26 : _GEN_384; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_386 = 5'h1b == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_27 : _GEN_385; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_387 = 5'h1c == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_28 : _GEN_386; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_388 = 5'h1d == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_29 : _GEN_387; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_389 = 5'h1e == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_30 : _GEN_388; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_20 = 5'h1f == _myTriMemVec2_20_T_1[4:0] ? myTriMemVec_31 : _GEN_389; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_19_T_1 = 16'hc + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_392 = 5'h1 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_393 = 5'h2 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_2 : _GEN_392; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_394 = 5'h3 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_3 : _GEN_393; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_395 = 5'h4 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_4 : _GEN_394; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_396 = 5'h5 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_5 : _GEN_395; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_397 = 5'h6 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_6 : _GEN_396; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_398 = 5'h7 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_7 : _GEN_397; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_399 = 5'h8 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_8 : _GEN_398; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_400 = 5'h9 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_9 : _GEN_399; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_401 = 5'ha == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_10 : _GEN_400; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_402 = 5'hb == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_11 : _GEN_401; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_403 = 5'hc == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_12 : _GEN_402; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_404 = 5'hd == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_13 : _GEN_403; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_405 = 5'he == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_14 : _GEN_404; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_406 = 5'hf == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_15 : _GEN_405; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_407 = 5'h10 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_16 : _GEN_406; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_408 = 5'h11 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_17 : _GEN_407; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_409 = 5'h12 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_18 : _GEN_408; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_410 = 5'h13 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_19 : _GEN_409; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_411 = 5'h14 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_20 : _GEN_410; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_412 = 5'h15 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_21 : _GEN_411; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_413 = 5'h16 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_22 : _GEN_412; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_414 = 5'h17 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_23 : _GEN_413; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_415 = 5'h18 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_24 : _GEN_414; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_416 = 5'h19 == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_25 : _GEN_415; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_417 = 5'h1a == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_26 : _GEN_416; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_418 = 5'h1b == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_27 : _GEN_417; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_419 = 5'h1c == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_28 : _GEN_418; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_420 = 5'h1d == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_29 : _GEN_419; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_421 = 5'h1e == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_30 : _GEN_420; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_19 = 5'h1f == _myTriMemVec2_19_T_1[4:0] ? myTriMemVec_31 : _GEN_421; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_18_T_1 = 16'hd + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_424 = 5'h1 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_425 = 5'h2 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_2 : _GEN_424; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_426 = 5'h3 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_3 : _GEN_425; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_427 = 5'h4 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_4 : _GEN_426; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_428 = 5'h5 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_5 : _GEN_427; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_429 = 5'h6 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_6 : _GEN_428; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_430 = 5'h7 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_7 : _GEN_429; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_431 = 5'h8 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_8 : _GEN_430; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_432 = 5'h9 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_9 : _GEN_431; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_433 = 5'ha == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_10 : _GEN_432; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_434 = 5'hb == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_11 : _GEN_433; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_435 = 5'hc == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_12 : _GEN_434; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_436 = 5'hd == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_13 : _GEN_435; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_437 = 5'he == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_14 : _GEN_436; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_438 = 5'hf == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_15 : _GEN_437; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_439 = 5'h10 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_16 : _GEN_438; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_440 = 5'h11 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_17 : _GEN_439; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_441 = 5'h12 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_18 : _GEN_440; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_442 = 5'h13 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_19 : _GEN_441; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_443 = 5'h14 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_20 : _GEN_442; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_444 = 5'h15 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_21 : _GEN_443; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_445 = 5'h16 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_22 : _GEN_444; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_446 = 5'h17 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_23 : _GEN_445; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_447 = 5'h18 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_24 : _GEN_446; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_448 = 5'h19 == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_25 : _GEN_447; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_449 = 5'h1a == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_26 : _GEN_448; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_450 = 5'h1b == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_27 : _GEN_449; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_451 = 5'h1c == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_28 : _GEN_450; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_452 = 5'h1d == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_29 : _GEN_451; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_453 = 5'h1e == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_30 : _GEN_452; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_18 = 5'h1f == _myTriMemVec2_18_T_1[4:0] ? myTriMemVec_31 : _GEN_453; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_17_T_1 = 16'he + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_456 = 5'h1 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_457 = 5'h2 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_2 : _GEN_456; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_458 = 5'h3 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_3 : _GEN_457; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_459 = 5'h4 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_4 : _GEN_458; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_460 = 5'h5 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_5 : _GEN_459; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_461 = 5'h6 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_6 : _GEN_460; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_462 = 5'h7 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_7 : _GEN_461; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_463 = 5'h8 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_8 : _GEN_462; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_464 = 5'h9 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_9 : _GEN_463; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_465 = 5'ha == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_10 : _GEN_464; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_466 = 5'hb == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_11 : _GEN_465; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_467 = 5'hc == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_12 : _GEN_466; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_468 = 5'hd == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_13 : _GEN_467; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_469 = 5'he == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_14 : _GEN_468; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_470 = 5'hf == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_15 : _GEN_469; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_471 = 5'h10 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_16 : _GEN_470; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_472 = 5'h11 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_17 : _GEN_471; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_473 = 5'h12 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_18 : _GEN_472; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_474 = 5'h13 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_19 : _GEN_473; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_475 = 5'h14 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_20 : _GEN_474; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_476 = 5'h15 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_21 : _GEN_475; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_477 = 5'h16 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_22 : _GEN_476; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_478 = 5'h17 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_23 : _GEN_477; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_479 = 5'h18 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_24 : _GEN_478; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_480 = 5'h19 == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_25 : _GEN_479; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_481 = 5'h1a == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_26 : _GEN_480; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_482 = 5'h1b == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_27 : _GEN_481; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_483 = 5'h1c == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_28 : _GEN_482; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_484 = 5'h1d == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_29 : _GEN_483; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_485 = 5'h1e == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_30 : _GEN_484; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_17 = 5'h1f == _myTriMemVec2_17_T_1[4:0] ? myTriMemVec_31 : _GEN_485; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_16_T_1 = 16'hf + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_488 = 5'h1 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_489 = 5'h2 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_2 : _GEN_488; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_490 = 5'h3 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_3 : _GEN_489; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_491 = 5'h4 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_4 : _GEN_490; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_492 = 5'h5 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_5 : _GEN_491; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_493 = 5'h6 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_6 : _GEN_492; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_494 = 5'h7 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_7 : _GEN_493; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_495 = 5'h8 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_8 : _GEN_494; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_496 = 5'h9 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_9 : _GEN_495; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_497 = 5'ha == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_10 : _GEN_496; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_498 = 5'hb == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_11 : _GEN_497; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_499 = 5'hc == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_12 : _GEN_498; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_500 = 5'hd == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_13 : _GEN_499; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_501 = 5'he == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_14 : _GEN_500; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_502 = 5'hf == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_15 : _GEN_501; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_503 = 5'h10 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_16 : _GEN_502; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_504 = 5'h11 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_17 : _GEN_503; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_505 = 5'h12 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_18 : _GEN_504; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_506 = 5'h13 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_19 : _GEN_505; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_507 = 5'h14 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_20 : _GEN_506; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_508 = 5'h15 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_21 : _GEN_507; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_509 = 5'h16 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_22 : _GEN_508; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_510 = 5'h17 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_23 : _GEN_509; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_511 = 5'h18 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_24 : _GEN_510; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_512 = 5'h19 == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_25 : _GEN_511; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_513 = 5'h1a == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_26 : _GEN_512; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_514 = 5'h1b == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_27 : _GEN_513; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_515 = 5'h1c == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_28 : _GEN_514; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_516 = 5'h1d == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_29 : _GEN_515; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_517 = 5'h1e == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_30 : _GEN_516; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_16 = 5'h1f == _myTriMemVec2_16_T_1[4:0] ? myTriMemVec_31 : _GEN_517; // @[hh_core.scala 127:{54,54}]
  wire [255:0] myTriMemWire_hi_lo = {myTriMemVec2_23,myTriMemVec2_22,myTriMemVec2_21,myTriMemVec2_20,myTriMemVec2_19,
    myTriMemVec2_18,myTriMemVec2_17,myTriMemVec2_16}; // @[hh_core.scala 131:42]
  wire [15:0] _myTriMemVec2_15_T_1 = 16'h10 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_520 = 5'h1 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_521 = 5'h2 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_2 : _GEN_520; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_522 = 5'h3 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_3 : _GEN_521; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_523 = 5'h4 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_4 : _GEN_522; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_524 = 5'h5 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_5 : _GEN_523; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_525 = 5'h6 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_6 : _GEN_524; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_526 = 5'h7 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_7 : _GEN_525; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_527 = 5'h8 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_8 : _GEN_526; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_528 = 5'h9 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_9 : _GEN_527; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_529 = 5'ha == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_10 : _GEN_528; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_530 = 5'hb == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_11 : _GEN_529; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_531 = 5'hc == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_12 : _GEN_530; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_532 = 5'hd == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_13 : _GEN_531; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_533 = 5'he == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_14 : _GEN_532; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_534 = 5'hf == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_15 : _GEN_533; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_535 = 5'h10 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_16 : _GEN_534; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_536 = 5'h11 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_17 : _GEN_535; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_537 = 5'h12 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_18 : _GEN_536; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_538 = 5'h13 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_19 : _GEN_537; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_539 = 5'h14 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_20 : _GEN_538; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_540 = 5'h15 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_21 : _GEN_539; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_541 = 5'h16 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_22 : _GEN_540; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_542 = 5'h17 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_23 : _GEN_541; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_543 = 5'h18 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_24 : _GEN_542; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_544 = 5'h19 == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_25 : _GEN_543; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_545 = 5'h1a == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_26 : _GEN_544; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_546 = 5'h1b == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_27 : _GEN_545; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_547 = 5'h1c == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_28 : _GEN_546; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_548 = 5'h1d == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_29 : _GEN_547; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_549 = 5'h1e == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_30 : _GEN_548; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_15 = 5'h1f == _myTriMemVec2_15_T_1[4:0] ? myTriMemVec_31 : _GEN_549; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_14_T_1 = 16'h11 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_552 = 5'h1 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_553 = 5'h2 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_2 : _GEN_552; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_554 = 5'h3 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_3 : _GEN_553; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_555 = 5'h4 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_4 : _GEN_554; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_556 = 5'h5 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_5 : _GEN_555; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_557 = 5'h6 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_6 : _GEN_556; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_558 = 5'h7 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_7 : _GEN_557; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_559 = 5'h8 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_8 : _GEN_558; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_560 = 5'h9 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_9 : _GEN_559; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_561 = 5'ha == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_10 : _GEN_560; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_562 = 5'hb == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_11 : _GEN_561; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_563 = 5'hc == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_12 : _GEN_562; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_564 = 5'hd == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_13 : _GEN_563; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_565 = 5'he == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_14 : _GEN_564; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_566 = 5'hf == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_15 : _GEN_565; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_567 = 5'h10 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_16 : _GEN_566; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_568 = 5'h11 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_17 : _GEN_567; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_569 = 5'h12 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_18 : _GEN_568; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_570 = 5'h13 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_19 : _GEN_569; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_571 = 5'h14 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_20 : _GEN_570; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_572 = 5'h15 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_21 : _GEN_571; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_573 = 5'h16 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_22 : _GEN_572; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_574 = 5'h17 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_23 : _GEN_573; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_575 = 5'h18 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_24 : _GEN_574; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_576 = 5'h19 == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_25 : _GEN_575; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_577 = 5'h1a == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_26 : _GEN_576; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_578 = 5'h1b == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_27 : _GEN_577; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_579 = 5'h1c == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_28 : _GEN_578; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_580 = 5'h1d == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_29 : _GEN_579; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_581 = 5'h1e == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_30 : _GEN_580; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_14 = 5'h1f == _myTriMemVec2_14_T_1[4:0] ? myTriMemVec_31 : _GEN_581; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_13_T_1 = 16'h12 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_584 = 5'h1 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_585 = 5'h2 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_2 : _GEN_584; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_586 = 5'h3 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_3 : _GEN_585; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_587 = 5'h4 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_4 : _GEN_586; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_588 = 5'h5 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_5 : _GEN_587; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_589 = 5'h6 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_6 : _GEN_588; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_590 = 5'h7 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_7 : _GEN_589; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_591 = 5'h8 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_8 : _GEN_590; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_592 = 5'h9 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_9 : _GEN_591; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_593 = 5'ha == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_10 : _GEN_592; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_594 = 5'hb == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_11 : _GEN_593; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_595 = 5'hc == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_12 : _GEN_594; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_596 = 5'hd == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_13 : _GEN_595; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_597 = 5'he == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_14 : _GEN_596; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_598 = 5'hf == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_15 : _GEN_597; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_599 = 5'h10 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_16 : _GEN_598; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_600 = 5'h11 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_17 : _GEN_599; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_601 = 5'h12 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_18 : _GEN_600; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_602 = 5'h13 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_19 : _GEN_601; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_603 = 5'h14 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_20 : _GEN_602; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_604 = 5'h15 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_21 : _GEN_603; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_605 = 5'h16 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_22 : _GEN_604; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_606 = 5'h17 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_23 : _GEN_605; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_607 = 5'h18 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_24 : _GEN_606; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_608 = 5'h19 == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_25 : _GEN_607; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_609 = 5'h1a == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_26 : _GEN_608; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_610 = 5'h1b == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_27 : _GEN_609; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_611 = 5'h1c == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_28 : _GEN_610; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_612 = 5'h1d == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_29 : _GEN_611; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_613 = 5'h1e == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_30 : _GEN_612; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_13 = 5'h1f == _myTriMemVec2_13_T_1[4:0] ? myTriMemVec_31 : _GEN_613; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_12_T_1 = 16'h13 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_616 = 5'h1 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_617 = 5'h2 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_2 : _GEN_616; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_618 = 5'h3 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_3 : _GEN_617; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_619 = 5'h4 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_4 : _GEN_618; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_620 = 5'h5 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_5 : _GEN_619; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_621 = 5'h6 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_6 : _GEN_620; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_622 = 5'h7 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_7 : _GEN_621; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_623 = 5'h8 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_8 : _GEN_622; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_624 = 5'h9 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_9 : _GEN_623; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_625 = 5'ha == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_10 : _GEN_624; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_626 = 5'hb == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_11 : _GEN_625; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_627 = 5'hc == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_12 : _GEN_626; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_628 = 5'hd == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_13 : _GEN_627; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_629 = 5'he == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_14 : _GEN_628; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_630 = 5'hf == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_15 : _GEN_629; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_631 = 5'h10 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_16 : _GEN_630; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_632 = 5'h11 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_17 : _GEN_631; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_633 = 5'h12 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_18 : _GEN_632; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_634 = 5'h13 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_19 : _GEN_633; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_635 = 5'h14 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_20 : _GEN_634; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_636 = 5'h15 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_21 : _GEN_635; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_637 = 5'h16 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_22 : _GEN_636; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_638 = 5'h17 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_23 : _GEN_637; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_639 = 5'h18 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_24 : _GEN_638; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_640 = 5'h19 == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_25 : _GEN_639; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_641 = 5'h1a == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_26 : _GEN_640; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_642 = 5'h1b == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_27 : _GEN_641; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_643 = 5'h1c == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_28 : _GEN_642; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_644 = 5'h1d == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_29 : _GEN_643; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_645 = 5'h1e == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_30 : _GEN_644; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_12 = 5'h1f == _myTriMemVec2_12_T_1[4:0] ? myTriMemVec_31 : _GEN_645; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_11_T_1 = 16'h14 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_648 = 5'h1 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_649 = 5'h2 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_2 : _GEN_648; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_650 = 5'h3 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_3 : _GEN_649; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_651 = 5'h4 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_4 : _GEN_650; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_652 = 5'h5 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_5 : _GEN_651; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_653 = 5'h6 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_6 : _GEN_652; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_654 = 5'h7 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_7 : _GEN_653; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_655 = 5'h8 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_8 : _GEN_654; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_656 = 5'h9 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_9 : _GEN_655; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_657 = 5'ha == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_10 : _GEN_656; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_658 = 5'hb == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_11 : _GEN_657; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_659 = 5'hc == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_12 : _GEN_658; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_660 = 5'hd == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_13 : _GEN_659; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_661 = 5'he == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_14 : _GEN_660; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_662 = 5'hf == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_15 : _GEN_661; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_663 = 5'h10 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_16 : _GEN_662; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_664 = 5'h11 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_17 : _GEN_663; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_665 = 5'h12 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_18 : _GEN_664; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_666 = 5'h13 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_19 : _GEN_665; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_667 = 5'h14 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_20 : _GEN_666; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_668 = 5'h15 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_21 : _GEN_667; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_669 = 5'h16 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_22 : _GEN_668; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_670 = 5'h17 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_23 : _GEN_669; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_671 = 5'h18 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_24 : _GEN_670; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_672 = 5'h19 == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_25 : _GEN_671; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_673 = 5'h1a == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_26 : _GEN_672; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_674 = 5'h1b == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_27 : _GEN_673; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_675 = 5'h1c == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_28 : _GEN_674; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_676 = 5'h1d == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_29 : _GEN_675; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_677 = 5'h1e == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_30 : _GEN_676; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_11 = 5'h1f == _myTriMemVec2_11_T_1[4:0] ? myTriMemVec_31 : _GEN_677; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_10_T_1 = 16'h15 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_680 = 5'h1 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_681 = 5'h2 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_2 : _GEN_680; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_682 = 5'h3 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_3 : _GEN_681; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_683 = 5'h4 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_4 : _GEN_682; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_684 = 5'h5 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_5 : _GEN_683; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_685 = 5'h6 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_6 : _GEN_684; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_686 = 5'h7 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_7 : _GEN_685; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_687 = 5'h8 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_8 : _GEN_686; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_688 = 5'h9 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_9 : _GEN_687; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_689 = 5'ha == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_10 : _GEN_688; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_690 = 5'hb == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_11 : _GEN_689; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_691 = 5'hc == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_12 : _GEN_690; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_692 = 5'hd == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_13 : _GEN_691; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_693 = 5'he == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_14 : _GEN_692; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_694 = 5'hf == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_15 : _GEN_693; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_695 = 5'h10 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_16 : _GEN_694; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_696 = 5'h11 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_17 : _GEN_695; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_697 = 5'h12 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_18 : _GEN_696; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_698 = 5'h13 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_19 : _GEN_697; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_699 = 5'h14 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_20 : _GEN_698; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_700 = 5'h15 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_21 : _GEN_699; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_701 = 5'h16 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_22 : _GEN_700; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_702 = 5'h17 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_23 : _GEN_701; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_703 = 5'h18 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_24 : _GEN_702; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_704 = 5'h19 == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_25 : _GEN_703; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_705 = 5'h1a == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_26 : _GEN_704; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_706 = 5'h1b == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_27 : _GEN_705; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_707 = 5'h1c == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_28 : _GEN_706; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_708 = 5'h1d == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_29 : _GEN_707; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_709 = 5'h1e == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_30 : _GEN_708; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_10 = 5'h1f == _myTriMemVec2_10_T_1[4:0] ? myTriMemVec_31 : _GEN_709; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_9_T_1 = 16'h16 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_712 = 5'h1 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_713 = 5'h2 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_2 : _GEN_712; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_714 = 5'h3 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_3 : _GEN_713; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_715 = 5'h4 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_4 : _GEN_714; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_716 = 5'h5 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_5 : _GEN_715; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_717 = 5'h6 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_6 : _GEN_716; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_718 = 5'h7 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_7 : _GEN_717; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_719 = 5'h8 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_8 : _GEN_718; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_720 = 5'h9 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_9 : _GEN_719; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_721 = 5'ha == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_10 : _GEN_720; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_722 = 5'hb == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_11 : _GEN_721; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_723 = 5'hc == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_12 : _GEN_722; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_724 = 5'hd == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_13 : _GEN_723; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_725 = 5'he == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_14 : _GEN_724; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_726 = 5'hf == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_15 : _GEN_725; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_727 = 5'h10 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_16 : _GEN_726; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_728 = 5'h11 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_17 : _GEN_727; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_729 = 5'h12 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_18 : _GEN_728; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_730 = 5'h13 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_19 : _GEN_729; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_731 = 5'h14 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_20 : _GEN_730; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_732 = 5'h15 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_21 : _GEN_731; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_733 = 5'h16 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_22 : _GEN_732; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_734 = 5'h17 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_23 : _GEN_733; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_735 = 5'h18 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_24 : _GEN_734; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_736 = 5'h19 == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_25 : _GEN_735; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_737 = 5'h1a == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_26 : _GEN_736; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_738 = 5'h1b == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_27 : _GEN_737; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_739 = 5'h1c == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_28 : _GEN_738; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_740 = 5'h1d == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_29 : _GEN_739; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_741 = 5'h1e == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_30 : _GEN_740; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_9 = 5'h1f == _myTriMemVec2_9_T_1[4:0] ? myTriMemVec_31 : _GEN_741; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_8_T_1 = 16'h17 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_744 = 5'h1 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_745 = 5'h2 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_2 : _GEN_744; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_746 = 5'h3 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_3 : _GEN_745; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_747 = 5'h4 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_4 : _GEN_746; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_748 = 5'h5 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_5 : _GEN_747; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_749 = 5'h6 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_6 : _GEN_748; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_750 = 5'h7 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_7 : _GEN_749; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_751 = 5'h8 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_8 : _GEN_750; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_752 = 5'h9 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_9 : _GEN_751; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_753 = 5'ha == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_10 : _GEN_752; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_754 = 5'hb == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_11 : _GEN_753; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_755 = 5'hc == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_12 : _GEN_754; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_756 = 5'hd == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_13 : _GEN_755; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_757 = 5'he == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_14 : _GEN_756; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_758 = 5'hf == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_15 : _GEN_757; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_759 = 5'h10 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_16 : _GEN_758; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_760 = 5'h11 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_17 : _GEN_759; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_761 = 5'h12 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_18 : _GEN_760; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_762 = 5'h13 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_19 : _GEN_761; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_763 = 5'h14 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_20 : _GEN_762; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_764 = 5'h15 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_21 : _GEN_763; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_765 = 5'h16 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_22 : _GEN_764; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_766 = 5'h17 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_23 : _GEN_765; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_767 = 5'h18 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_24 : _GEN_766; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_768 = 5'h19 == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_25 : _GEN_767; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_769 = 5'h1a == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_26 : _GEN_768; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_770 = 5'h1b == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_27 : _GEN_769; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_771 = 5'h1c == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_28 : _GEN_770; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_772 = 5'h1d == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_29 : _GEN_771; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_773 = 5'h1e == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_30 : _GEN_772; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_8 = 5'h1f == _myTriMemVec2_8_T_1[4:0] ? myTriMemVec_31 : _GEN_773; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_7_T_1 = 16'h18 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_776 = 5'h1 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_777 = 5'h2 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_2 : _GEN_776; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_778 = 5'h3 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_3 : _GEN_777; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_779 = 5'h4 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_4 : _GEN_778; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_780 = 5'h5 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_5 : _GEN_779; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_781 = 5'h6 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_6 : _GEN_780; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_782 = 5'h7 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_7 : _GEN_781; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_783 = 5'h8 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_8 : _GEN_782; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_784 = 5'h9 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_9 : _GEN_783; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_785 = 5'ha == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_10 : _GEN_784; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_786 = 5'hb == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_11 : _GEN_785; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_787 = 5'hc == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_12 : _GEN_786; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_788 = 5'hd == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_13 : _GEN_787; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_789 = 5'he == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_14 : _GEN_788; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_790 = 5'hf == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_15 : _GEN_789; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_791 = 5'h10 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_16 : _GEN_790; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_792 = 5'h11 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_17 : _GEN_791; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_793 = 5'h12 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_18 : _GEN_792; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_794 = 5'h13 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_19 : _GEN_793; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_795 = 5'h14 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_20 : _GEN_794; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_796 = 5'h15 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_21 : _GEN_795; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_797 = 5'h16 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_22 : _GEN_796; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_798 = 5'h17 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_23 : _GEN_797; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_799 = 5'h18 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_24 : _GEN_798; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_800 = 5'h19 == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_25 : _GEN_799; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_801 = 5'h1a == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_26 : _GEN_800; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_802 = 5'h1b == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_27 : _GEN_801; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_803 = 5'h1c == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_28 : _GEN_802; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_804 = 5'h1d == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_29 : _GEN_803; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_805 = 5'h1e == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_30 : _GEN_804; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_7 = 5'h1f == _myTriMemVec2_7_T_1[4:0] ? myTriMemVec_31 : _GEN_805; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_6_T_1 = 16'h19 + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_808 = 5'h1 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_809 = 5'h2 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_2 : _GEN_808; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_810 = 5'h3 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_3 : _GEN_809; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_811 = 5'h4 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_4 : _GEN_810; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_812 = 5'h5 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_5 : _GEN_811; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_813 = 5'h6 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_6 : _GEN_812; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_814 = 5'h7 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_7 : _GEN_813; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_815 = 5'h8 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_8 : _GEN_814; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_816 = 5'h9 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_9 : _GEN_815; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_817 = 5'ha == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_10 : _GEN_816; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_818 = 5'hb == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_11 : _GEN_817; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_819 = 5'hc == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_12 : _GEN_818; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_820 = 5'hd == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_13 : _GEN_819; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_821 = 5'he == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_14 : _GEN_820; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_822 = 5'hf == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_15 : _GEN_821; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_823 = 5'h10 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_16 : _GEN_822; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_824 = 5'h11 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_17 : _GEN_823; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_825 = 5'h12 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_18 : _GEN_824; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_826 = 5'h13 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_19 : _GEN_825; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_827 = 5'h14 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_20 : _GEN_826; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_828 = 5'h15 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_21 : _GEN_827; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_829 = 5'h16 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_22 : _GEN_828; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_830 = 5'h17 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_23 : _GEN_829; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_831 = 5'h18 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_24 : _GEN_830; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_832 = 5'h19 == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_25 : _GEN_831; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_833 = 5'h1a == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_26 : _GEN_832; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_834 = 5'h1b == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_27 : _GEN_833; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_835 = 5'h1c == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_28 : _GEN_834; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_836 = 5'h1d == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_29 : _GEN_835; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_837 = 5'h1e == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_30 : _GEN_836; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_6 = 5'h1f == _myTriMemVec2_6_T_1[4:0] ? myTriMemVec_31 : _GEN_837; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_5_T_1 = 16'h1a + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_840 = 5'h1 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_841 = 5'h2 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_2 : _GEN_840; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_842 = 5'h3 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_3 : _GEN_841; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_843 = 5'h4 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_4 : _GEN_842; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_844 = 5'h5 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_5 : _GEN_843; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_845 = 5'h6 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_6 : _GEN_844; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_846 = 5'h7 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_7 : _GEN_845; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_847 = 5'h8 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_8 : _GEN_846; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_848 = 5'h9 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_9 : _GEN_847; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_849 = 5'ha == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_10 : _GEN_848; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_850 = 5'hb == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_11 : _GEN_849; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_851 = 5'hc == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_12 : _GEN_850; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_852 = 5'hd == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_13 : _GEN_851; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_853 = 5'he == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_14 : _GEN_852; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_854 = 5'hf == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_15 : _GEN_853; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_855 = 5'h10 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_16 : _GEN_854; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_856 = 5'h11 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_17 : _GEN_855; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_857 = 5'h12 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_18 : _GEN_856; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_858 = 5'h13 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_19 : _GEN_857; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_859 = 5'h14 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_20 : _GEN_858; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_860 = 5'h15 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_21 : _GEN_859; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_861 = 5'h16 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_22 : _GEN_860; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_862 = 5'h17 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_23 : _GEN_861; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_863 = 5'h18 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_24 : _GEN_862; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_864 = 5'h19 == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_25 : _GEN_863; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_865 = 5'h1a == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_26 : _GEN_864; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_866 = 5'h1b == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_27 : _GEN_865; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_867 = 5'h1c == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_28 : _GEN_866; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_868 = 5'h1d == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_29 : _GEN_867; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_869 = 5'h1e == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_30 : _GEN_868; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_5 = 5'h1f == _myTriMemVec2_5_T_1[4:0] ? myTriMemVec_31 : _GEN_869; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_4_T_1 = 16'h1b + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_872 = 5'h1 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_873 = 5'h2 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_2 : _GEN_872; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_874 = 5'h3 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_3 : _GEN_873; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_875 = 5'h4 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_4 : _GEN_874; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_876 = 5'h5 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_5 : _GEN_875; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_877 = 5'h6 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_6 : _GEN_876; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_878 = 5'h7 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_7 : _GEN_877; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_879 = 5'h8 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_8 : _GEN_878; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_880 = 5'h9 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_9 : _GEN_879; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_881 = 5'ha == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_10 : _GEN_880; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_882 = 5'hb == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_11 : _GEN_881; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_883 = 5'hc == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_12 : _GEN_882; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_884 = 5'hd == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_13 : _GEN_883; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_885 = 5'he == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_14 : _GEN_884; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_886 = 5'hf == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_15 : _GEN_885; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_887 = 5'h10 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_16 : _GEN_886; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_888 = 5'h11 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_17 : _GEN_887; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_889 = 5'h12 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_18 : _GEN_888; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_890 = 5'h13 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_19 : _GEN_889; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_891 = 5'h14 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_20 : _GEN_890; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_892 = 5'h15 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_21 : _GEN_891; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_893 = 5'h16 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_22 : _GEN_892; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_894 = 5'h17 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_23 : _GEN_893; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_895 = 5'h18 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_24 : _GEN_894; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_896 = 5'h19 == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_25 : _GEN_895; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_897 = 5'h1a == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_26 : _GEN_896; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_898 = 5'h1b == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_27 : _GEN_897; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_899 = 5'h1c == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_28 : _GEN_898; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_900 = 5'h1d == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_29 : _GEN_899; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_901 = 5'h1e == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_30 : _GEN_900; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_4 = 5'h1f == _myTriMemVec2_4_T_1[4:0] ? myTriMemVec_31 : _GEN_901; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_3_T_1 = 16'h1c + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_904 = 5'h1 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_905 = 5'h2 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_2 : _GEN_904; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_906 = 5'h3 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_3 : _GEN_905; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_907 = 5'h4 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_4 : _GEN_906; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_908 = 5'h5 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_5 : _GEN_907; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_909 = 5'h6 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_6 : _GEN_908; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_910 = 5'h7 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_7 : _GEN_909; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_911 = 5'h8 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_8 : _GEN_910; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_912 = 5'h9 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_9 : _GEN_911; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_913 = 5'ha == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_10 : _GEN_912; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_914 = 5'hb == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_11 : _GEN_913; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_915 = 5'hc == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_12 : _GEN_914; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_916 = 5'hd == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_13 : _GEN_915; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_917 = 5'he == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_14 : _GEN_916; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_918 = 5'hf == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_15 : _GEN_917; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_919 = 5'h10 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_16 : _GEN_918; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_920 = 5'h11 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_17 : _GEN_919; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_921 = 5'h12 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_18 : _GEN_920; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_922 = 5'h13 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_19 : _GEN_921; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_923 = 5'h14 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_20 : _GEN_922; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_924 = 5'h15 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_21 : _GEN_923; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_925 = 5'h16 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_22 : _GEN_924; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_926 = 5'h17 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_23 : _GEN_925; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_927 = 5'h18 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_24 : _GEN_926; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_928 = 5'h19 == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_25 : _GEN_927; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_929 = 5'h1a == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_26 : _GEN_928; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_930 = 5'h1b == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_27 : _GEN_929; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_931 = 5'h1c == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_28 : _GEN_930; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_932 = 5'h1d == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_29 : _GEN_931; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_933 = 5'h1e == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_30 : _GEN_932; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_3 = 5'h1f == _myTriMemVec2_3_T_1[4:0] ? myTriMemVec_31 : _GEN_933; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_2_T_1 = 16'h1d + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_936 = 5'h1 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_937 = 5'h2 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_2 : _GEN_936; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_938 = 5'h3 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_3 : _GEN_937; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_939 = 5'h4 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_4 : _GEN_938; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_940 = 5'h5 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_5 : _GEN_939; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_941 = 5'h6 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_6 : _GEN_940; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_942 = 5'h7 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_7 : _GEN_941; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_943 = 5'h8 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_8 : _GEN_942; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_944 = 5'h9 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_9 : _GEN_943; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_945 = 5'ha == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_10 : _GEN_944; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_946 = 5'hb == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_11 : _GEN_945; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_947 = 5'hc == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_12 : _GEN_946; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_948 = 5'hd == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_13 : _GEN_947; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_949 = 5'he == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_14 : _GEN_948; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_950 = 5'hf == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_15 : _GEN_949; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_951 = 5'h10 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_16 : _GEN_950; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_952 = 5'h11 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_17 : _GEN_951; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_953 = 5'h12 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_18 : _GEN_952; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_954 = 5'h13 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_19 : _GEN_953; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_955 = 5'h14 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_20 : _GEN_954; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_956 = 5'h15 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_21 : _GEN_955; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_957 = 5'h16 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_22 : _GEN_956; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_958 = 5'h17 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_23 : _GEN_957; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_959 = 5'h18 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_24 : _GEN_958; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_960 = 5'h19 == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_25 : _GEN_959; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_961 = 5'h1a == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_26 : _GEN_960; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_962 = 5'h1b == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_27 : _GEN_961; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_963 = 5'h1c == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_28 : _GEN_962; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_964 = 5'h1d == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_29 : _GEN_963; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_965 = 5'h1e == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_30 : _GEN_964; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_2 = 5'h1f == _myTriMemVec2_2_T_1[4:0] ? myTriMemVec_31 : _GEN_965; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_1_T_1 = 16'h1e + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_968 = 5'h1 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_969 = 5'h2 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_2 : _GEN_968; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_970 = 5'h3 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_3 : _GEN_969; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_971 = 5'h4 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_4 : _GEN_970; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_972 = 5'h5 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_5 : _GEN_971; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_973 = 5'h6 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_6 : _GEN_972; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_974 = 5'h7 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_7 : _GEN_973; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_975 = 5'h8 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_8 : _GEN_974; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_976 = 5'h9 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_9 : _GEN_975; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_977 = 5'ha == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_10 : _GEN_976; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_978 = 5'hb == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_11 : _GEN_977; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_979 = 5'hc == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_12 : _GEN_978; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_980 = 5'hd == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_13 : _GEN_979; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_981 = 5'he == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_14 : _GEN_980; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_982 = 5'hf == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_15 : _GEN_981; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_983 = 5'h10 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_16 : _GEN_982; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_984 = 5'h11 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_17 : _GEN_983; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_985 = 5'h12 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_18 : _GEN_984; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_986 = 5'h13 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_19 : _GEN_985; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_987 = 5'h14 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_20 : _GEN_986; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_988 = 5'h15 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_21 : _GEN_987; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_989 = 5'h16 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_22 : _GEN_988; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_990 = 5'h17 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_23 : _GEN_989; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_991 = 5'h18 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_24 : _GEN_990; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_992 = 5'h19 == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_25 : _GEN_991; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_993 = 5'h1a == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_26 : _GEN_992; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_994 = 5'h1b == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_27 : _GEN_993; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_995 = 5'h1c == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_28 : _GEN_994; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_996 = 5'h1d == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_29 : _GEN_995; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_997 = 5'h1e == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_30 : _GEN_996; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_1 = 5'h1f == _myTriMemVec2_1_T_1[4:0] ? myTriMemVec_31 : _GEN_997; // @[hh_core.scala 127:{54,54}]
  wire [15:0] _myTriMemVec2_0_T_1 = 16'h1f + io_hh_cnt; // @[hh_core.scala 127:74]
  wire [31:0] _GEN_1000 = 5'h1 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_1 : myTriMemVec_0; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1001 = 5'h2 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_2 : _GEN_1000; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1002 = 5'h3 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_3 : _GEN_1001; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1003 = 5'h4 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_4 : _GEN_1002; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1004 = 5'h5 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_5 : _GEN_1003; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1005 = 5'h6 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_6 : _GEN_1004; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1006 = 5'h7 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_7 : _GEN_1005; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1007 = 5'h8 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_8 : _GEN_1006; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1008 = 5'h9 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_9 : _GEN_1007; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1009 = 5'ha == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_10 : _GEN_1008; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1010 = 5'hb == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_11 : _GEN_1009; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1011 = 5'hc == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_12 : _GEN_1010; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1012 = 5'hd == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_13 : _GEN_1011; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1013 = 5'he == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_14 : _GEN_1012; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1014 = 5'hf == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_15 : _GEN_1013; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1015 = 5'h10 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_16 : _GEN_1014; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1016 = 5'h11 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_17 : _GEN_1015; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1017 = 5'h12 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_18 : _GEN_1016; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1018 = 5'h13 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_19 : _GEN_1017; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1019 = 5'h14 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_20 : _GEN_1018; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1020 = 5'h15 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_21 : _GEN_1019; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1021 = 5'h16 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_22 : _GEN_1020; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1022 = 5'h17 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_23 : _GEN_1021; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1023 = 5'h18 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_24 : _GEN_1022; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1024 = 5'h19 == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_25 : _GEN_1023; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1025 = 5'h1a == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_26 : _GEN_1024; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1026 = 5'h1b == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_27 : _GEN_1025; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1027 = 5'h1c == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_28 : _GEN_1026; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1028 = 5'h1d == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_29 : _GEN_1027; // @[hh_core.scala 127:{54,54}]
  wire [31:0] _GEN_1029 = 5'h1e == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_30 : _GEN_1028; // @[hh_core.scala 127:{54,54}]
  wire [31:0] myTriMemVec2_0 = 5'h1f == _myTriMemVec2_0_T_1[4:0] ? myTriMemVec_31 : _GEN_1029; // @[hh_core.scala 127:{54,54}]
  wire [255:0] myTriMemWire_lo_lo = {myTriMemVec2_7,myTriMemVec2_6,myTriMemVec2_5,myTriMemVec2_4,myTriMemVec2_3,
    myTriMemVec2_2,myTriMemVec2_1,myTriMemVec2_0}; // @[hh_core.scala 131:42]
  wire [511:0] myTriMemWire_lo = {myTriMemVec2_15,myTriMemVec2_14,myTriMemVec2_13,myTriMemVec2_12,myTriMemVec2_11,
    myTriMemVec2_10,myTriMemVec2_9,myTriMemVec2_8,myTriMemWire_lo_lo}; // @[hh_core.scala 131:42]
  wire [1023:0] myTriMemWire = {myTriMemVec2_31,myTriMemVec2_30,myTriMemVec2_29,myTriMemVec2_28,myTriMemVec2_27,
    myTriMemVec2_26,myTriMemVec2_25,myTriMemVec2_24,myTriMemWire_hi_lo,myTriMemWire_lo}; // @[hh_core.scala 131:42]
  wire [21:0] _hh_din_update_T = io_hh_cnt * 6'h20; // @[hh_core.scala 134:65]
  wire [1023:0] _hh_din_update_T_1 = myTriMemWire >> _hh_din_update_T; // @[hh_core.scala 134:52]
  wire [1023:0] _GEN_5 = hh1_din_rdy ? io_dmx1_mem_doutb : 1024'h0; // @[hh_core.scala 113:36 114:31 116:31]
  wire [1023:0] dmx_mem_doutb = hh0_din_rdy ? io_dmx0_mem_doutb : _GEN_5; // @[hh_core.scala 111:30 112:31]
  wire [2047:0] _hh_din_update_T_2 = {_hh_din_update_T_1,dmx_mem_doutb}; // @[Cat.scala 31:58]
  wire [31:0] myHhdoutVec_63 = io_hh_dout[31:0]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_62 = io_hh_dout[63:32]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_61 = io_hh_dout[95:64]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_60 = io_hh_dout[127:96]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_59 = io_hh_dout[159:128]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_58 = io_hh_dout[191:160]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_57 = io_hh_dout[223:192]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_56 = io_hh_dout[255:224]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_55 = io_hh_dout[287:256]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_54 = io_hh_dout[319:288]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_53 = io_hh_dout[351:320]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_52 = io_hh_dout[383:352]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_51 = io_hh_dout[415:384]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_50 = io_hh_dout[447:416]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_49 = io_hh_dout[479:448]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_48 = io_hh_dout[511:480]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_47 = io_hh_dout[543:512]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_46 = io_hh_dout[575:544]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_45 = io_hh_dout[607:576]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_44 = io_hh_dout[639:608]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_43 = io_hh_dout[671:640]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_42 = io_hh_dout[703:672]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_41 = io_hh_dout[735:704]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_40 = io_hh_dout[767:736]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_39 = io_hh_dout[799:768]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_38 = io_hh_dout[831:800]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_37 = io_hh_dout[863:832]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_36 = io_hh_dout[895:864]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_35 = io_hh_dout[927:896]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_34 = io_hh_dout[959:928]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_33 = io_hh_dout[991:960]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_32 = io_hh_dout[1023:992]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_31 = io_hh_dout[1055:1024]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_30 = io_hh_dout[1087:1056]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_29 = io_hh_dout[1119:1088]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_28 = io_hh_dout[1151:1120]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_27 = io_hh_dout[1183:1152]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_26 = io_hh_dout[1215:1184]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_25 = io_hh_dout[1247:1216]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_24 = io_hh_dout[1279:1248]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_23 = io_hh_dout[1311:1280]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_22 = io_hh_dout[1343:1312]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_21 = io_hh_dout[1375:1344]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_20 = io_hh_dout[1407:1376]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_19 = io_hh_dout[1439:1408]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_18 = io_hh_dout[1471:1440]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_17 = io_hh_dout[1503:1472]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_16 = io_hh_dout[1535:1504]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_15 = io_hh_dout[1567:1536]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_14 = io_hh_dout[1599:1568]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_13 = io_hh_dout[1631:1600]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_12 = io_hh_dout[1663:1632]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_11 = io_hh_dout[1695:1664]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_10 = io_hh_dout[1727:1696]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_9 = io_hh_dout[1759:1728]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_8 = io_hh_dout[1791:1760]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_7 = io_hh_dout[1823:1792]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_6 = io_hh_dout[1855:1824]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_5 = io_hh_dout[1887:1856]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_4 = io_hh_dout[1919:1888]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_3 = io_hh_dout[1951:1920]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_2 = io_hh_dout[1983:1952]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_1 = io_hh_dout[2015:1984]; // @[hh_core.scala 144:45]
  wire [31:0] myHhdoutVec_0 = io_hh_dout[2047:2016]; // @[hh_core.scala 144:45]
  wire [31:0] _GEN_1034 = 6'h1 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1035 = 6'h2 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_2 : _GEN_1034; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1036 = 6'h3 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_3 : _GEN_1035; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1037 = 6'h4 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_4 : _GEN_1036; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1038 = 6'h5 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_5 : _GEN_1037; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1039 = 6'h6 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_6 : _GEN_1038; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1040 = 6'h7 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_7 : _GEN_1039; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1041 = 6'h8 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_8 : _GEN_1040; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1042 = 6'h9 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_9 : _GEN_1041; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1043 = 6'ha == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_10 : _GEN_1042; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1044 = 6'hb == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_11 : _GEN_1043; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1045 = 6'hc == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_12 : _GEN_1044; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1046 = 6'hd == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_13 : _GEN_1045; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1047 = 6'he == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_14 : _GEN_1046; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1048 = 6'hf == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_15 : _GEN_1047; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1049 = 6'h10 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_16 : _GEN_1048; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1050 = 6'h11 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_17 : _GEN_1049; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1051 = 6'h12 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_18 : _GEN_1050; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1052 = 6'h13 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_19 : _GEN_1051; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1053 = 6'h14 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_20 : _GEN_1052; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1054 = 6'h15 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_21 : _GEN_1053; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1055 = 6'h16 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_22 : _GEN_1054; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1056 = 6'h17 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_23 : _GEN_1055; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1057 = 6'h18 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_24 : _GEN_1056; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1058 = 6'h19 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_25 : _GEN_1057; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1059 = 6'h1a == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_26 : _GEN_1058; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1060 = 6'h1b == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_27 : _GEN_1059; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1061 = 6'h1c == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_28 : _GEN_1060; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1062 = 6'h1d == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_29 : _GEN_1061; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1063 = 6'h1e == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_30 : _GEN_1062; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1064 = 6'h1f == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_31 : _GEN_1063; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1065 = 6'h20 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_32 : _GEN_1064; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1066 = 6'h21 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_33 : _GEN_1065; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1067 = 6'h22 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_34 : _GEN_1066; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1068 = 6'h23 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_35 : _GEN_1067; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1069 = 6'h24 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_36 : _GEN_1068; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1070 = 6'h25 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_37 : _GEN_1069; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1071 = 6'h26 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_38 : _GEN_1070; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1072 = 6'h27 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_39 : _GEN_1071; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1073 = 6'h28 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_40 : _GEN_1072; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1074 = 6'h29 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_41 : _GEN_1073; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1075 = 6'h2a == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_42 : _GEN_1074; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1076 = 6'h2b == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_43 : _GEN_1075; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1077 = 6'h2c == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_44 : _GEN_1076; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1078 = 6'h2d == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_45 : _GEN_1077; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1079 = 6'h2e == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_46 : _GEN_1078; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1080 = 6'h2f == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_47 : _GEN_1079; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1081 = 6'h30 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_48 : _GEN_1080; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1082 = 6'h31 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_49 : _GEN_1081; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1083 = 6'h32 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_50 : _GEN_1082; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1084 = 6'h33 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_51 : _GEN_1083; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1085 = 6'h34 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_52 : _GEN_1084; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1086 = 6'h35 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_53 : _GEN_1085; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1087 = 6'h36 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_54 : _GEN_1086; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1088 = 6'h37 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_55 : _GEN_1087; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1089 = 6'h38 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_56 : _GEN_1088; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1090 = 6'h39 == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_57 : _GEN_1089; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1091 = 6'h3a == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_58 : _GEN_1090; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1092 = 6'h3b == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_59 : _GEN_1091; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1093 = 6'h3c == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_60 : _GEN_1092; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1094 = 6'h3d == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_61 : _GEN_1093; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1095 = 6'h3e == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_62 : _GEN_1094; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_63 = 6'h3f == _myTriMemVec2_31_T[5:0] ? myHhdoutVec_63 : _GEN_1095; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1098 = 6'h1 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1099 = 6'h2 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_2 : _GEN_1098; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1100 = 6'h3 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_3 : _GEN_1099; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1101 = 6'h4 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_4 : _GEN_1100; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1102 = 6'h5 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_5 : _GEN_1101; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1103 = 6'h6 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_6 : _GEN_1102; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1104 = 6'h7 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_7 : _GEN_1103; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1105 = 6'h8 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_8 : _GEN_1104; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1106 = 6'h9 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_9 : _GEN_1105; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1107 = 6'ha == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_10 : _GEN_1106; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1108 = 6'hb == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_11 : _GEN_1107; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1109 = 6'hc == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_12 : _GEN_1108; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1110 = 6'hd == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_13 : _GEN_1109; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1111 = 6'he == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_14 : _GEN_1110; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1112 = 6'hf == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_15 : _GEN_1111; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1113 = 6'h10 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_16 : _GEN_1112; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1114 = 6'h11 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_17 : _GEN_1113; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1115 = 6'h12 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_18 : _GEN_1114; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1116 = 6'h13 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_19 : _GEN_1115; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1117 = 6'h14 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_20 : _GEN_1116; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1118 = 6'h15 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_21 : _GEN_1117; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1119 = 6'h16 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_22 : _GEN_1118; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1120 = 6'h17 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_23 : _GEN_1119; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1121 = 6'h18 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_24 : _GEN_1120; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1122 = 6'h19 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_25 : _GEN_1121; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1123 = 6'h1a == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_26 : _GEN_1122; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1124 = 6'h1b == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_27 : _GEN_1123; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1125 = 6'h1c == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_28 : _GEN_1124; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1126 = 6'h1d == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_29 : _GEN_1125; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1127 = 6'h1e == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_30 : _GEN_1126; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1128 = 6'h1f == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_31 : _GEN_1127; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1129 = 6'h20 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_32 : _GEN_1128; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1130 = 6'h21 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_33 : _GEN_1129; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1131 = 6'h22 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_34 : _GEN_1130; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1132 = 6'h23 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_35 : _GEN_1131; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1133 = 6'h24 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_36 : _GEN_1132; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1134 = 6'h25 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_37 : _GEN_1133; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1135 = 6'h26 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_38 : _GEN_1134; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1136 = 6'h27 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_39 : _GEN_1135; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1137 = 6'h28 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_40 : _GEN_1136; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1138 = 6'h29 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_41 : _GEN_1137; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1139 = 6'h2a == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_42 : _GEN_1138; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1140 = 6'h2b == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_43 : _GEN_1139; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1141 = 6'h2c == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_44 : _GEN_1140; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1142 = 6'h2d == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_45 : _GEN_1141; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1143 = 6'h2e == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_46 : _GEN_1142; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1144 = 6'h2f == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_47 : _GEN_1143; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1145 = 6'h30 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_48 : _GEN_1144; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1146 = 6'h31 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_49 : _GEN_1145; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1147 = 6'h32 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_50 : _GEN_1146; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1148 = 6'h33 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_51 : _GEN_1147; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1149 = 6'h34 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_52 : _GEN_1148; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1150 = 6'h35 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_53 : _GEN_1149; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1151 = 6'h36 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_54 : _GEN_1150; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1152 = 6'h37 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_55 : _GEN_1151; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1153 = 6'h38 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_56 : _GEN_1152; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1154 = 6'h39 == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_57 : _GEN_1153; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1155 = 6'h3a == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_58 : _GEN_1154; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1156 = 6'h3b == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_59 : _GEN_1155; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1157 = 6'h3c == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_60 : _GEN_1156; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1158 = 6'h3d == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_61 : _GEN_1157; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1159 = 6'h3e == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_62 : _GEN_1158; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_62 = 6'h3f == _myTriMemVec2_30_T_1[5:0] ? myHhdoutVec_63 : _GEN_1159; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1162 = 6'h1 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1163 = 6'h2 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_2 : _GEN_1162; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1164 = 6'h3 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_3 : _GEN_1163; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1165 = 6'h4 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_4 : _GEN_1164; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1166 = 6'h5 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_5 : _GEN_1165; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1167 = 6'h6 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_6 : _GEN_1166; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1168 = 6'h7 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_7 : _GEN_1167; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1169 = 6'h8 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_8 : _GEN_1168; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1170 = 6'h9 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_9 : _GEN_1169; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1171 = 6'ha == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_10 : _GEN_1170; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1172 = 6'hb == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_11 : _GEN_1171; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1173 = 6'hc == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_12 : _GEN_1172; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1174 = 6'hd == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_13 : _GEN_1173; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1175 = 6'he == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_14 : _GEN_1174; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1176 = 6'hf == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_15 : _GEN_1175; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1177 = 6'h10 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_16 : _GEN_1176; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1178 = 6'h11 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_17 : _GEN_1177; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1179 = 6'h12 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_18 : _GEN_1178; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1180 = 6'h13 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_19 : _GEN_1179; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1181 = 6'h14 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_20 : _GEN_1180; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1182 = 6'h15 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_21 : _GEN_1181; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1183 = 6'h16 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_22 : _GEN_1182; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1184 = 6'h17 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_23 : _GEN_1183; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1185 = 6'h18 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_24 : _GEN_1184; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1186 = 6'h19 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_25 : _GEN_1185; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1187 = 6'h1a == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_26 : _GEN_1186; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1188 = 6'h1b == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_27 : _GEN_1187; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1189 = 6'h1c == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_28 : _GEN_1188; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1190 = 6'h1d == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_29 : _GEN_1189; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1191 = 6'h1e == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_30 : _GEN_1190; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1192 = 6'h1f == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_31 : _GEN_1191; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1193 = 6'h20 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_32 : _GEN_1192; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1194 = 6'h21 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_33 : _GEN_1193; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1195 = 6'h22 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_34 : _GEN_1194; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1196 = 6'h23 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_35 : _GEN_1195; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1197 = 6'h24 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_36 : _GEN_1196; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1198 = 6'h25 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_37 : _GEN_1197; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1199 = 6'h26 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_38 : _GEN_1198; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1200 = 6'h27 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_39 : _GEN_1199; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1201 = 6'h28 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_40 : _GEN_1200; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1202 = 6'h29 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_41 : _GEN_1201; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1203 = 6'h2a == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_42 : _GEN_1202; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1204 = 6'h2b == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_43 : _GEN_1203; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1205 = 6'h2c == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_44 : _GEN_1204; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1206 = 6'h2d == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_45 : _GEN_1205; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1207 = 6'h2e == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_46 : _GEN_1206; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1208 = 6'h2f == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_47 : _GEN_1207; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1209 = 6'h30 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_48 : _GEN_1208; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1210 = 6'h31 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_49 : _GEN_1209; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1211 = 6'h32 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_50 : _GEN_1210; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1212 = 6'h33 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_51 : _GEN_1211; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1213 = 6'h34 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_52 : _GEN_1212; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1214 = 6'h35 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_53 : _GEN_1213; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1215 = 6'h36 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_54 : _GEN_1214; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1216 = 6'h37 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_55 : _GEN_1215; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1217 = 6'h38 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_56 : _GEN_1216; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1218 = 6'h39 == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_57 : _GEN_1217; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1219 = 6'h3a == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_58 : _GEN_1218; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1220 = 6'h3b == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_59 : _GEN_1219; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1221 = 6'h3c == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_60 : _GEN_1220; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1222 = 6'h3d == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_61 : _GEN_1221; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1223 = 6'h3e == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_62 : _GEN_1222; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_61 = 6'h3f == _myTriMemVec2_29_T_1[5:0] ? myHhdoutVec_63 : _GEN_1223; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1226 = 6'h1 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1227 = 6'h2 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_2 : _GEN_1226; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1228 = 6'h3 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_3 : _GEN_1227; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1229 = 6'h4 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_4 : _GEN_1228; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1230 = 6'h5 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_5 : _GEN_1229; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1231 = 6'h6 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_6 : _GEN_1230; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1232 = 6'h7 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_7 : _GEN_1231; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1233 = 6'h8 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_8 : _GEN_1232; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1234 = 6'h9 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_9 : _GEN_1233; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1235 = 6'ha == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_10 : _GEN_1234; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1236 = 6'hb == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_11 : _GEN_1235; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1237 = 6'hc == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_12 : _GEN_1236; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1238 = 6'hd == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_13 : _GEN_1237; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1239 = 6'he == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_14 : _GEN_1238; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1240 = 6'hf == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_15 : _GEN_1239; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1241 = 6'h10 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_16 : _GEN_1240; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1242 = 6'h11 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_17 : _GEN_1241; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1243 = 6'h12 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_18 : _GEN_1242; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1244 = 6'h13 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_19 : _GEN_1243; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1245 = 6'h14 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_20 : _GEN_1244; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1246 = 6'h15 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_21 : _GEN_1245; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1247 = 6'h16 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_22 : _GEN_1246; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1248 = 6'h17 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_23 : _GEN_1247; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1249 = 6'h18 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_24 : _GEN_1248; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1250 = 6'h19 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_25 : _GEN_1249; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1251 = 6'h1a == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_26 : _GEN_1250; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1252 = 6'h1b == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_27 : _GEN_1251; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1253 = 6'h1c == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_28 : _GEN_1252; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1254 = 6'h1d == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_29 : _GEN_1253; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1255 = 6'h1e == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_30 : _GEN_1254; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1256 = 6'h1f == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_31 : _GEN_1255; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1257 = 6'h20 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_32 : _GEN_1256; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1258 = 6'h21 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_33 : _GEN_1257; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1259 = 6'h22 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_34 : _GEN_1258; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1260 = 6'h23 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_35 : _GEN_1259; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1261 = 6'h24 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_36 : _GEN_1260; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1262 = 6'h25 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_37 : _GEN_1261; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1263 = 6'h26 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_38 : _GEN_1262; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1264 = 6'h27 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_39 : _GEN_1263; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1265 = 6'h28 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_40 : _GEN_1264; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1266 = 6'h29 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_41 : _GEN_1265; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1267 = 6'h2a == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_42 : _GEN_1266; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1268 = 6'h2b == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_43 : _GEN_1267; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1269 = 6'h2c == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_44 : _GEN_1268; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1270 = 6'h2d == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_45 : _GEN_1269; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1271 = 6'h2e == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_46 : _GEN_1270; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1272 = 6'h2f == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_47 : _GEN_1271; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1273 = 6'h30 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_48 : _GEN_1272; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1274 = 6'h31 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_49 : _GEN_1273; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1275 = 6'h32 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_50 : _GEN_1274; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1276 = 6'h33 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_51 : _GEN_1275; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1277 = 6'h34 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_52 : _GEN_1276; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1278 = 6'h35 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_53 : _GEN_1277; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1279 = 6'h36 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_54 : _GEN_1278; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1280 = 6'h37 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_55 : _GEN_1279; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1281 = 6'h38 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_56 : _GEN_1280; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1282 = 6'h39 == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_57 : _GEN_1281; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1283 = 6'h3a == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_58 : _GEN_1282; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1284 = 6'h3b == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_59 : _GEN_1283; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1285 = 6'h3c == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_60 : _GEN_1284; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1286 = 6'h3d == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_61 : _GEN_1285; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1287 = 6'h3e == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_62 : _GEN_1286; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_60 = 6'h3f == _myTriMemVec2_28_T_1[5:0] ? myHhdoutVec_63 : _GEN_1287; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1290 = 6'h1 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1291 = 6'h2 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_2 : _GEN_1290; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1292 = 6'h3 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_3 : _GEN_1291; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1293 = 6'h4 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_4 : _GEN_1292; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1294 = 6'h5 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_5 : _GEN_1293; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1295 = 6'h6 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_6 : _GEN_1294; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1296 = 6'h7 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_7 : _GEN_1295; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1297 = 6'h8 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_8 : _GEN_1296; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1298 = 6'h9 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_9 : _GEN_1297; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1299 = 6'ha == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_10 : _GEN_1298; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1300 = 6'hb == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_11 : _GEN_1299; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1301 = 6'hc == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_12 : _GEN_1300; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1302 = 6'hd == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_13 : _GEN_1301; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1303 = 6'he == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_14 : _GEN_1302; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1304 = 6'hf == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_15 : _GEN_1303; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1305 = 6'h10 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_16 : _GEN_1304; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1306 = 6'h11 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_17 : _GEN_1305; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1307 = 6'h12 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_18 : _GEN_1306; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1308 = 6'h13 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_19 : _GEN_1307; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1309 = 6'h14 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_20 : _GEN_1308; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1310 = 6'h15 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_21 : _GEN_1309; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1311 = 6'h16 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_22 : _GEN_1310; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1312 = 6'h17 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_23 : _GEN_1311; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1313 = 6'h18 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_24 : _GEN_1312; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1314 = 6'h19 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_25 : _GEN_1313; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1315 = 6'h1a == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_26 : _GEN_1314; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1316 = 6'h1b == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_27 : _GEN_1315; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1317 = 6'h1c == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_28 : _GEN_1316; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1318 = 6'h1d == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_29 : _GEN_1317; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1319 = 6'h1e == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_30 : _GEN_1318; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1320 = 6'h1f == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_31 : _GEN_1319; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1321 = 6'h20 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_32 : _GEN_1320; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1322 = 6'h21 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_33 : _GEN_1321; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1323 = 6'h22 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_34 : _GEN_1322; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1324 = 6'h23 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_35 : _GEN_1323; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1325 = 6'h24 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_36 : _GEN_1324; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1326 = 6'h25 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_37 : _GEN_1325; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1327 = 6'h26 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_38 : _GEN_1326; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1328 = 6'h27 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_39 : _GEN_1327; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1329 = 6'h28 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_40 : _GEN_1328; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1330 = 6'h29 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_41 : _GEN_1329; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1331 = 6'h2a == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_42 : _GEN_1330; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1332 = 6'h2b == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_43 : _GEN_1331; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1333 = 6'h2c == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_44 : _GEN_1332; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1334 = 6'h2d == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_45 : _GEN_1333; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1335 = 6'h2e == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_46 : _GEN_1334; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1336 = 6'h2f == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_47 : _GEN_1335; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1337 = 6'h30 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_48 : _GEN_1336; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1338 = 6'h31 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_49 : _GEN_1337; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1339 = 6'h32 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_50 : _GEN_1338; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1340 = 6'h33 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_51 : _GEN_1339; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1341 = 6'h34 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_52 : _GEN_1340; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1342 = 6'h35 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_53 : _GEN_1341; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1343 = 6'h36 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_54 : _GEN_1342; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1344 = 6'h37 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_55 : _GEN_1343; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1345 = 6'h38 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_56 : _GEN_1344; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1346 = 6'h39 == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_57 : _GEN_1345; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1347 = 6'h3a == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_58 : _GEN_1346; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1348 = 6'h3b == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_59 : _GEN_1347; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1349 = 6'h3c == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_60 : _GEN_1348; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1350 = 6'h3d == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_61 : _GEN_1349; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1351 = 6'h3e == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_62 : _GEN_1350; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_59 = 6'h3f == _myTriMemVec2_27_T_1[5:0] ? myHhdoutVec_63 : _GEN_1351; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1354 = 6'h1 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1355 = 6'h2 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_2 : _GEN_1354; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1356 = 6'h3 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_3 : _GEN_1355; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1357 = 6'h4 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_4 : _GEN_1356; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1358 = 6'h5 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_5 : _GEN_1357; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1359 = 6'h6 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_6 : _GEN_1358; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1360 = 6'h7 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_7 : _GEN_1359; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1361 = 6'h8 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_8 : _GEN_1360; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1362 = 6'h9 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_9 : _GEN_1361; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1363 = 6'ha == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_10 : _GEN_1362; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1364 = 6'hb == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_11 : _GEN_1363; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1365 = 6'hc == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_12 : _GEN_1364; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1366 = 6'hd == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_13 : _GEN_1365; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1367 = 6'he == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_14 : _GEN_1366; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1368 = 6'hf == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_15 : _GEN_1367; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1369 = 6'h10 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_16 : _GEN_1368; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1370 = 6'h11 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_17 : _GEN_1369; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1371 = 6'h12 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_18 : _GEN_1370; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1372 = 6'h13 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_19 : _GEN_1371; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1373 = 6'h14 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_20 : _GEN_1372; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1374 = 6'h15 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_21 : _GEN_1373; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1375 = 6'h16 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_22 : _GEN_1374; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1376 = 6'h17 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_23 : _GEN_1375; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1377 = 6'h18 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_24 : _GEN_1376; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1378 = 6'h19 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_25 : _GEN_1377; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1379 = 6'h1a == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_26 : _GEN_1378; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1380 = 6'h1b == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_27 : _GEN_1379; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1381 = 6'h1c == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_28 : _GEN_1380; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1382 = 6'h1d == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_29 : _GEN_1381; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1383 = 6'h1e == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_30 : _GEN_1382; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1384 = 6'h1f == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_31 : _GEN_1383; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1385 = 6'h20 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_32 : _GEN_1384; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1386 = 6'h21 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_33 : _GEN_1385; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1387 = 6'h22 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_34 : _GEN_1386; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1388 = 6'h23 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_35 : _GEN_1387; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1389 = 6'h24 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_36 : _GEN_1388; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1390 = 6'h25 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_37 : _GEN_1389; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1391 = 6'h26 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_38 : _GEN_1390; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1392 = 6'h27 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_39 : _GEN_1391; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1393 = 6'h28 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_40 : _GEN_1392; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1394 = 6'h29 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_41 : _GEN_1393; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1395 = 6'h2a == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_42 : _GEN_1394; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1396 = 6'h2b == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_43 : _GEN_1395; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1397 = 6'h2c == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_44 : _GEN_1396; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1398 = 6'h2d == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_45 : _GEN_1397; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1399 = 6'h2e == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_46 : _GEN_1398; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1400 = 6'h2f == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_47 : _GEN_1399; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1401 = 6'h30 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_48 : _GEN_1400; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1402 = 6'h31 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_49 : _GEN_1401; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1403 = 6'h32 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_50 : _GEN_1402; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1404 = 6'h33 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_51 : _GEN_1403; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1405 = 6'h34 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_52 : _GEN_1404; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1406 = 6'h35 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_53 : _GEN_1405; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1407 = 6'h36 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_54 : _GEN_1406; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1408 = 6'h37 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_55 : _GEN_1407; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1409 = 6'h38 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_56 : _GEN_1408; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1410 = 6'h39 == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_57 : _GEN_1409; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1411 = 6'h3a == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_58 : _GEN_1410; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1412 = 6'h3b == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_59 : _GEN_1411; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1413 = 6'h3c == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_60 : _GEN_1412; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1414 = 6'h3d == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_61 : _GEN_1413; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1415 = 6'h3e == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_62 : _GEN_1414; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_58 = 6'h3f == _myTriMemVec2_26_T_1[5:0] ? myHhdoutVec_63 : _GEN_1415; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1418 = 6'h1 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1419 = 6'h2 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_2 : _GEN_1418; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1420 = 6'h3 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_3 : _GEN_1419; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1421 = 6'h4 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_4 : _GEN_1420; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1422 = 6'h5 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_5 : _GEN_1421; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1423 = 6'h6 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_6 : _GEN_1422; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1424 = 6'h7 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_7 : _GEN_1423; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1425 = 6'h8 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_8 : _GEN_1424; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1426 = 6'h9 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_9 : _GEN_1425; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1427 = 6'ha == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_10 : _GEN_1426; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1428 = 6'hb == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_11 : _GEN_1427; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1429 = 6'hc == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_12 : _GEN_1428; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1430 = 6'hd == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_13 : _GEN_1429; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1431 = 6'he == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_14 : _GEN_1430; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1432 = 6'hf == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_15 : _GEN_1431; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1433 = 6'h10 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_16 : _GEN_1432; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1434 = 6'h11 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_17 : _GEN_1433; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1435 = 6'h12 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_18 : _GEN_1434; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1436 = 6'h13 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_19 : _GEN_1435; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1437 = 6'h14 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_20 : _GEN_1436; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1438 = 6'h15 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_21 : _GEN_1437; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1439 = 6'h16 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_22 : _GEN_1438; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1440 = 6'h17 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_23 : _GEN_1439; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1441 = 6'h18 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_24 : _GEN_1440; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1442 = 6'h19 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_25 : _GEN_1441; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1443 = 6'h1a == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_26 : _GEN_1442; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1444 = 6'h1b == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_27 : _GEN_1443; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1445 = 6'h1c == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_28 : _GEN_1444; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1446 = 6'h1d == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_29 : _GEN_1445; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1447 = 6'h1e == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_30 : _GEN_1446; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1448 = 6'h1f == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_31 : _GEN_1447; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1449 = 6'h20 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_32 : _GEN_1448; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1450 = 6'h21 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_33 : _GEN_1449; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1451 = 6'h22 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_34 : _GEN_1450; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1452 = 6'h23 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_35 : _GEN_1451; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1453 = 6'h24 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_36 : _GEN_1452; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1454 = 6'h25 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_37 : _GEN_1453; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1455 = 6'h26 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_38 : _GEN_1454; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1456 = 6'h27 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_39 : _GEN_1455; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1457 = 6'h28 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_40 : _GEN_1456; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1458 = 6'h29 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_41 : _GEN_1457; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1459 = 6'h2a == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_42 : _GEN_1458; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1460 = 6'h2b == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_43 : _GEN_1459; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1461 = 6'h2c == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_44 : _GEN_1460; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1462 = 6'h2d == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_45 : _GEN_1461; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1463 = 6'h2e == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_46 : _GEN_1462; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1464 = 6'h2f == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_47 : _GEN_1463; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1465 = 6'h30 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_48 : _GEN_1464; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1466 = 6'h31 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_49 : _GEN_1465; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1467 = 6'h32 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_50 : _GEN_1466; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1468 = 6'h33 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_51 : _GEN_1467; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1469 = 6'h34 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_52 : _GEN_1468; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1470 = 6'h35 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_53 : _GEN_1469; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1471 = 6'h36 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_54 : _GEN_1470; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1472 = 6'h37 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_55 : _GEN_1471; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1473 = 6'h38 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_56 : _GEN_1472; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1474 = 6'h39 == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_57 : _GEN_1473; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1475 = 6'h3a == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_58 : _GEN_1474; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1476 = 6'h3b == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_59 : _GEN_1475; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1477 = 6'h3c == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_60 : _GEN_1476; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1478 = 6'h3d == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_61 : _GEN_1477; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1479 = 6'h3e == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_62 : _GEN_1478; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_57 = 6'h3f == _myTriMemVec2_25_T_1[5:0] ? myHhdoutVec_63 : _GEN_1479; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1482 = 6'h1 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1483 = 6'h2 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_2 : _GEN_1482; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1484 = 6'h3 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_3 : _GEN_1483; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1485 = 6'h4 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_4 : _GEN_1484; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1486 = 6'h5 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_5 : _GEN_1485; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1487 = 6'h6 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_6 : _GEN_1486; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1488 = 6'h7 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_7 : _GEN_1487; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1489 = 6'h8 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_8 : _GEN_1488; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1490 = 6'h9 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_9 : _GEN_1489; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1491 = 6'ha == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_10 : _GEN_1490; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1492 = 6'hb == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_11 : _GEN_1491; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1493 = 6'hc == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_12 : _GEN_1492; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1494 = 6'hd == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_13 : _GEN_1493; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1495 = 6'he == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_14 : _GEN_1494; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1496 = 6'hf == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_15 : _GEN_1495; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1497 = 6'h10 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_16 : _GEN_1496; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1498 = 6'h11 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_17 : _GEN_1497; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1499 = 6'h12 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_18 : _GEN_1498; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1500 = 6'h13 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_19 : _GEN_1499; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1501 = 6'h14 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_20 : _GEN_1500; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1502 = 6'h15 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_21 : _GEN_1501; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1503 = 6'h16 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_22 : _GEN_1502; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1504 = 6'h17 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_23 : _GEN_1503; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1505 = 6'h18 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_24 : _GEN_1504; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1506 = 6'h19 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_25 : _GEN_1505; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1507 = 6'h1a == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_26 : _GEN_1506; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1508 = 6'h1b == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_27 : _GEN_1507; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1509 = 6'h1c == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_28 : _GEN_1508; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1510 = 6'h1d == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_29 : _GEN_1509; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1511 = 6'h1e == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_30 : _GEN_1510; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1512 = 6'h1f == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_31 : _GEN_1511; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1513 = 6'h20 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_32 : _GEN_1512; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1514 = 6'h21 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_33 : _GEN_1513; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1515 = 6'h22 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_34 : _GEN_1514; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1516 = 6'h23 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_35 : _GEN_1515; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1517 = 6'h24 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_36 : _GEN_1516; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1518 = 6'h25 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_37 : _GEN_1517; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1519 = 6'h26 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_38 : _GEN_1518; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1520 = 6'h27 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_39 : _GEN_1519; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1521 = 6'h28 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_40 : _GEN_1520; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1522 = 6'h29 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_41 : _GEN_1521; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1523 = 6'h2a == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_42 : _GEN_1522; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1524 = 6'h2b == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_43 : _GEN_1523; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1525 = 6'h2c == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_44 : _GEN_1524; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1526 = 6'h2d == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_45 : _GEN_1525; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1527 = 6'h2e == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_46 : _GEN_1526; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1528 = 6'h2f == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_47 : _GEN_1527; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1529 = 6'h30 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_48 : _GEN_1528; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1530 = 6'h31 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_49 : _GEN_1529; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1531 = 6'h32 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_50 : _GEN_1530; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1532 = 6'h33 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_51 : _GEN_1531; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1533 = 6'h34 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_52 : _GEN_1532; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1534 = 6'h35 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_53 : _GEN_1533; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1535 = 6'h36 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_54 : _GEN_1534; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1536 = 6'h37 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_55 : _GEN_1535; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1537 = 6'h38 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_56 : _GEN_1536; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1538 = 6'h39 == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_57 : _GEN_1537; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1539 = 6'h3a == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_58 : _GEN_1538; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1540 = 6'h3b == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_59 : _GEN_1539; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1541 = 6'h3c == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_60 : _GEN_1540; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1542 = 6'h3d == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_61 : _GEN_1541; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1543 = 6'h3e == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_62 : _GEN_1542; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_56 = 6'h3f == _myTriMemVec2_24_T_1[5:0] ? myHhdoutVec_63 : _GEN_1543; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1546 = 6'h1 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1547 = 6'h2 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_2 : _GEN_1546; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1548 = 6'h3 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_3 : _GEN_1547; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1549 = 6'h4 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_4 : _GEN_1548; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1550 = 6'h5 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_5 : _GEN_1549; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1551 = 6'h6 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_6 : _GEN_1550; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1552 = 6'h7 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_7 : _GEN_1551; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1553 = 6'h8 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_8 : _GEN_1552; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1554 = 6'h9 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_9 : _GEN_1553; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1555 = 6'ha == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_10 : _GEN_1554; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1556 = 6'hb == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_11 : _GEN_1555; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1557 = 6'hc == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_12 : _GEN_1556; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1558 = 6'hd == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_13 : _GEN_1557; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1559 = 6'he == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_14 : _GEN_1558; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1560 = 6'hf == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_15 : _GEN_1559; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1561 = 6'h10 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_16 : _GEN_1560; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1562 = 6'h11 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_17 : _GEN_1561; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1563 = 6'h12 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_18 : _GEN_1562; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1564 = 6'h13 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_19 : _GEN_1563; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1565 = 6'h14 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_20 : _GEN_1564; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1566 = 6'h15 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_21 : _GEN_1565; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1567 = 6'h16 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_22 : _GEN_1566; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1568 = 6'h17 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_23 : _GEN_1567; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1569 = 6'h18 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_24 : _GEN_1568; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1570 = 6'h19 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_25 : _GEN_1569; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1571 = 6'h1a == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_26 : _GEN_1570; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1572 = 6'h1b == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_27 : _GEN_1571; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1573 = 6'h1c == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_28 : _GEN_1572; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1574 = 6'h1d == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_29 : _GEN_1573; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1575 = 6'h1e == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_30 : _GEN_1574; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1576 = 6'h1f == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_31 : _GEN_1575; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1577 = 6'h20 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_32 : _GEN_1576; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1578 = 6'h21 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_33 : _GEN_1577; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1579 = 6'h22 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_34 : _GEN_1578; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1580 = 6'h23 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_35 : _GEN_1579; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1581 = 6'h24 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_36 : _GEN_1580; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1582 = 6'h25 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_37 : _GEN_1581; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1583 = 6'h26 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_38 : _GEN_1582; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1584 = 6'h27 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_39 : _GEN_1583; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1585 = 6'h28 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_40 : _GEN_1584; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1586 = 6'h29 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_41 : _GEN_1585; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1587 = 6'h2a == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_42 : _GEN_1586; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1588 = 6'h2b == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_43 : _GEN_1587; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1589 = 6'h2c == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_44 : _GEN_1588; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1590 = 6'h2d == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_45 : _GEN_1589; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1591 = 6'h2e == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_46 : _GEN_1590; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1592 = 6'h2f == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_47 : _GEN_1591; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1593 = 6'h30 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_48 : _GEN_1592; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1594 = 6'h31 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_49 : _GEN_1593; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1595 = 6'h32 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_50 : _GEN_1594; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1596 = 6'h33 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_51 : _GEN_1595; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1597 = 6'h34 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_52 : _GEN_1596; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1598 = 6'h35 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_53 : _GEN_1597; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1599 = 6'h36 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_54 : _GEN_1598; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1600 = 6'h37 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_55 : _GEN_1599; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1601 = 6'h38 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_56 : _GEN_1600; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1602 = 6'h39 == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_57 : _GEN_1601; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1603 = 6'h3a == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_58 : _GEN_1602; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1604 = 6'h3b == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_59 : _GEN_1603; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1605 = 6'h3c == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_60 : _GEN_1604; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1606 = 6'h3d == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_61 : _GEN_1605; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1607 = 6'h3e == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_62 : _GEN_1606; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_55 = 6'h3f == _myTriMemVec2_23_T_1[5:0] ? myHhdoutVec_63 : _GEN_1607; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1610 = 6'h1 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1611 = 6'h2 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_2 : _GEN_1610; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1612 = 6'h3 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_3 : _GEN_1611; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1613 = 6'h4 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_4 : _GEN_1612; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1614 = 6'h5 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_5 : _GEN_1613; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1615 = 6'h6 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_6 : _GEN_1614; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1616 = 6'h7 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_7 : _GEN_1615; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1617 = 6'h8 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_8 : _GEN_1616; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1618 = 6'h9 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_9 : _GEN_1617; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1619 = 6'ha == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_10 : _GEN_1618; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1620 = 6'hb == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_11 : _GEN_1619; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1621 = 6'hc == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_12 : _GEN_1620; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1622 = 6'hd == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_13 : _GEN_1621; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1623 = 6'he == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_14 : _GEN_1622; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1624 = 6'hf == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_15 : _GEN_1623; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1625 = 6'h10 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_16 : _GEN_1624; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1626 = 6'h11 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_17 : _GEN_1625; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1627 = 6'h12 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_18 : _GEN_1626; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1628 = 6'h13 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_19 : _GEN_1627; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1629 = 6'h14 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_20 : _GEN_1628; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1630 = 6'h15 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_21 : _GEN_1629; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1631 = 6'h16 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_22 : _GEN_1630; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1632 = 6'h17 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_23 : _GEN_1631; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1633 = 6'h18 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_24 : _GEN_1632; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1634 = 6'h19 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_25 : _GEN_1633; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1635 = 6'h1a == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_26 : _GEN_1634; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1636 = 6'h1b == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_27 : _GEN_1635; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1637 = 6'h1c == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_28 : _GEN_1636; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1638 = 6'h1d == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_29 : _GEN_1637; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1639 = 6'h1e == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_30 : _GEN_1638; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1640 = 6'h1f == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_31 : _GEN_1639; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1641 = 6'h20 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_32 : _GEN_1640; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1642 = 6'h21 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_33 : _GEN_1641; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1643 = 6'h22 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_34 : _GEN_1642; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1644 = 6'h23 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_35 : _GEN_1643; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1645 = 6'h24 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_36 : _GEN_1644; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1646 = 6'h25 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_37 : _GEN_1645; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1647 = 6'h26 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_38 : _GEN_1646; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1648 = 6'h27 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_39 : _GEN_1647; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1649 = 6'h28 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_40 : _GEN_1648; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1650 = 6'h29 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_41 : _GEN_1649; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1651 = 6'h2a == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_42 : _GEN_1650; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1652 = 6'h2b == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_43 : _GEN_1651; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1653 = 6'h2c == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_44 : _GEN_1652; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1654 = 6'h2d == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_45 : _GEN_1653; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1655 = 6'h2e == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_46 : _GEN_1654; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1656 = 6'h2f == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_47 : _GEN_1655; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1657 = 6'h30 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_48 : _GEN_1656; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1658 = 6'h31 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_49 : _GEN_1657; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1659 = 6'h32 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_50 : _GEN_1658; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1660 = 6'h33 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_51 : _GEN_1659; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1661 = 6'h34 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_52 : _GEN_1660; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1662 = 6'h35 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_53 : _GEN_1661; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1663 = 6'h36 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_54 : _GEN_1662; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1664 = 6'h37 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_55 : _GEN_1663; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1665 = 6'h38 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_56 : _GEN_1664; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1666 = 6'h39 == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_57 : _GEN_1665; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1667 = 6'h3a == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_58 : _GEN_1666; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1668 = 6'h3b == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_59 : _GEN_1667; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1669 = 6'h3c == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_60 : _GEN_1668; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1670 = 6'h3d == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_61 : _GEN_1669; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1671 = 6'h3e == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_62 : _GEN_1670; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_54 = 6'h3f == _myTriMemVec2_22_T_1[5:0] ? myHhdoutVec_63 : _GEN_1671; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1674 = 6'h1 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1675 = 6'h2 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_2 : _GEN_1674; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1676 = 6'h3 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_3 : _GEN_1675; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1677 = 6'h4 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_4 : _GEN_1676; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1678 = 6'h5 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_5 : _GEN_1677; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1679 = 6'h6 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_6 : _GEN_1678; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1680 = 6'h7 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_7 : _GEN_1679; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1681 = 6'h8 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_8 : _GEN_1680; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1682 = 6'h9 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_9 : _GEN_1681; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1683 = 6'ha == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_10 : _GEN_1682; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1684 = 6'hb == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_11 : _GEN_1683; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1685 = 6'hc == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_12 : _GEN_1684; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1686 = 6'hd == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_13 : _GEN_1685; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1687 = 6'he == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_14 : _GEN_1686; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1688 = 6'hf == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_15 : _GEN_1687; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1689 = 6'h10 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_16 : _GEN_1688; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1690 = 6'h11 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_17 : _GEN_1689; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1691 = 6'h12 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_18 : _GEN_1690; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1692 = 6'h13 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_19 : _GEN_1691; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1693 = 6'h14 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_20 : _GEN_1692; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1694 = 6'h15 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_21 : _GEN_1693; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1695 = 6'h16 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_22 : _GEN_1694; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1696 = 6'h17 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_23 : _GEN_1695; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1697 = 6'h18 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_24 : _GEN_1696; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1698 = 6'h19 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_25 : _GEN_1697; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1699 = 6'h1a == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_26 : _GEN_1698; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1700 = 6'h1b == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_27 : _GEN_1699; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1701 = 6'h1c == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_28 : _GEN_1700; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1702 = 6'h1d == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_29 : _GEN_1701; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1703 = 6'h1e == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_30 : _GEN_1702; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1704 = 6'h1f == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_31 : _GEN_1703; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1705 = 6'h20 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_32 : _GEN_1704; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1706 = 6'h21 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_33 : _GEN_1705; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1707 = 6'h22 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_34 : _GEN_1706; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1708 = 6'h23 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_35 : _GEN_1707; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1709 = 6'h24 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_36 : _GEN_1708; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1710 = 6'h25 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_37 : _GEN_1709; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1711 = 6'h26 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_38 : _GEN_1710; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1712 = 6'h27 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_39 : _GEN_1711; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1713 = 6'h28 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_40 : _GEN_1712; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1714 = 6'h29 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_41 : _GEN_1713; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1715 = 6'h2a == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_42 : _GEN_1714; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1716 = 6'h2b == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_43 : _GEN_1715; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1717 = 6'h2c == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_44 : _GEN_1716; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1718 = 6'h2d == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_45 : _GEN_1717; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1719 = 6'h2e == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_46 : _GEN_1718; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1720 = 6'h2f == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_47 : _GEN_1719; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1721 = 6'h30 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_48 : _GEN_1720; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1722 = 6'h31 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_49 : _GEN_1721; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1723 = 6'h32 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_50 : _GEN_1722; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1724 = 6'h33 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_51 : _GEN_1723; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1725 = 6'h34 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_52 : _GEN_1724; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1726 = 6'h35 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_53 : _GEN_1725; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1727 = 6'h36 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_54 : _GEN_1726; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1728 = 6'h37 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_55 : _GEN_1727; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1729 = 6'h38 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_56 : _GEN_1728; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1730 = 6'h39 == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_57 : _GEN_1729; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1731 = 6'h3a == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_58 : _GEN_1730; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1732 = 6'h3b == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_59 : _GEN_1731; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1733 = 6'h3c == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_60 : _GEN_1732; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1734 = 6'h3d == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_61 : _GEN_1733; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1735 = 6'h3e == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_62 : _GEN_1734; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_53 = 6'h3f == _myTriMemVec2_21_T_1[5:0] ? myHhdoutVec_63 : _GEN_1735; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1738 = 6'h1 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1739 = 6'h2 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_2 : _GEN_1738; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1740 = 6'h3 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_3 : _GEN_1739; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1741 = 6'h4 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_4 : _GEN_1740; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1742 = 6'h5 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_5 : _GEN_1741; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1743 = 6'h6 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_6 : _GEN_1742; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1744 = 6'h7 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_7 : _GEN_1743; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1745 = 6'h8 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_8 : _GEN_1744; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1746 = 6'h9 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_9 : _GEN_1745; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1747 = 6'ha == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_10 : _GEN_1746; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1748 = 6'hb == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_11 : _GEN_1747; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1749 = 6'hc == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_12 : _GEN_1748; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1750 = 6'hd == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_13 : _GEN_1749; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1751 = 6'he == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_14 : _GEN_1750; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1752 = 6'hf == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_15 : _GEN_1751; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1753 = 6'h10 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_16 : _GEN_1752; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1754 = 6'h11 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_17 : _GEN_1753; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1755 = 6'h12 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_18 : _GEN_1754; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1756 = 6'h13 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_19 : _GEN_1755; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1757 = 6'h14 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_20 : _GEN_1756; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1758 = 6'h15 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_21 : _GEN_1757; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1759 = 6'h16 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_22 : _GEN_1758; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1760 = 6'h17 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_23 : _GEN_1759; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1761 = 6'h18 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_24 : _GEN_1760; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1762 = 6'h19 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_25 : _GEN_1761; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1763 = 6'h1a == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_26 : _GEN_1762; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1764 = 6'h1b == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_27 : _GEN_1763; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1765 = 6'h1c == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_28 : _GEN_1764; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1766 = 6'h1d == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_29 : _GEN_1765; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1767 = 6'h1e == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_30 : _GEN_1766; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1768 = 6'h1f == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_31 : _GEN_1767; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1769 = 6'h20 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_32 : _GEN_1768; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1770 = 6'h21 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_33 : _GEN_1769; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1771 = 6'h22 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_34 : _GEN_1770; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1772 = 6'h23 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_35 : _GEN_1771; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1773 = 6'h24 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_36 : _GEN_1772; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1774 = 6'h25 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_37 : _GEN_1773; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1775 = 6'h26 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_38 : _GEN_1774; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1776 = 6'h27 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_39 : _GEN_1775; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1777 = 6'h28 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_40 : _GEN_1776; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1778 = 6'h29 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_41 : _GEN_1777; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1779 = 6'h2a == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_42 : _GEN_1778; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1780 = 6'h2b == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_43 : _GEN_1779; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1781 = 6'h2c == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_44 : _GEN_1780; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1782 = 6'h2d == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_45 : _GEN_1781; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1783 = 6'h2e == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_46 : _GEN_1782; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1784 = 6'h2f == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_47 : _GEN_1783; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1785 = 6'h30 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_48 : _GEN_1784; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1786 = 6'h31 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_49 : _GEN_1785; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1787 = 6'h32 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_50 : _GEN_1786; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1788 = 6'h33 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_51 : _GEN_1787; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1789 = 6'h34 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_52 : _GEN_1788; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1790 = 6'h35 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_53 : _GEN_1789; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1791 = 6'h36 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_54 : _GEN_1790; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1792 = 6'h37 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_55 : _GEN_1791; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1793 = 6'h38 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_56 : _GEN_1792; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1794 = 6'h39 == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_57 : _GEN_1793; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1795 = 6'h3a == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_58 : _GEN_1794; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1796 = 6'h3b == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_59 : _GEN_1795; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1797 = 6'h3c == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_60 : _GEN_1796; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1798 = 6'h3d == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_61 : _GEN_1797; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1799 = 6'h3e == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_62 : _GEN_1798; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_52 = 6'h3f == _myTriMemVec2_20_T_1[5:0] ? myHhdoutVec_63 : _GEN_1799; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1802 = 6'h1 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1803 = 6'h2 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_2 : _GEN_1802; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1804 = 6'h3 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_3 : _GEN_1803; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1805 = 6'h4 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_4 : _GEN_1804; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1806 = 6'h5 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_5 : _GEN_1805; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1807 = 6'h6 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_6 : _GEN_1806; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1808 = 6'h7 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_7 : _GEN_1807; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1809 = 6'h8 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_8 : _GEN_1808; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1810 = 6'h9 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_9 : _GEN_1809; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1811 = 6'ha == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_10 : _GEN_1810; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1812 = 6'hb == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_11 : _GEN_1811; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1813 = 6'hc == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_12 : _GEN_1812; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1814 = 6'hd == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_13 : _GEN_1813; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1815 = 6'he == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_14 : _GEN_1814; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1816 = 6'hf == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_15 : _GEN_1815; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1817 = 6'h10 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_16 : _GEN_1816; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1818 = 6'h11 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_17 : _GEN_1817; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1819 = 6'h12 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_18 : _GEN_1818; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1820 = 6'h13 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_19 : _GEN_1819; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1821 = 6'h14 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_20 : _GEN_1820; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1822 = 6'h15 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_21 : _GEN_1821; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1823 = 6'h16 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_22 : _GEN_1822; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1824 = 6'h17 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_23 : _GEN_1823; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1825 = 6'h18 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_24 : _GEN_1824; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1826 = 6'h19 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_25 : _GEN_1825; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1827 = 6'h1a == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_26 : _GEN_1826; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1828 = 6'h1b == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_27 : _GEN_1827; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1829 = 6'h1c == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_28 : _GEN_1828; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1830 = 6'h1d == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_29 : _GEN_1829; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1831 = 6'h1e == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_30 : _GEN_1830; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1832 = 6'h1f == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_31 : _GEN_1831; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1833 = 6'h20 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_32 : _GEN_1832; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1834 = 6'h21 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_33 : _GEN_1833; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1835 = 6'h22 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_34 : _GEN_1834; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1836 = 6'h23 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_35 : _GEN_1835; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1837 = 6'h24 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_36 : _GEN_1836; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1838 = 6'h25 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_37 : _GEN_1837; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1839 = 6'h26 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_38 : _GEN_1838; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1840 = 6'h27 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_39 : _GEN_1839; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1841 = 6'h28 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_40 : _GEN_1840; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1842 = 6'h29 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_41 : _GEN_1841; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1843 = 6'h2a == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_42 : _GEN_1842; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1844 = 6'h2b == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_43 : _GEN_1843; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1845 = 6'h2c == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_44 : _GEN_1844; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1846 = 6'h2d == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_45 : _GEN_1845; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1847 = 6'h2e == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_46 : _GEN_1846; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1848 = 6'h2f == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_47 : _GEN_1847; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1849 = 6'h30 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_48 : _GEN_1848; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1850 = 6'h31 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_49 : _GEN_1849; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1851 = 6'h32 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_50 : _GEN_1850; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1852 = 6'h33 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_51 : _GEN_1851; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1853 = 6'h34 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_52 : _GEN_1852; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1854 = 6'h35 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_53 : _GEN_1853; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1855 = 6'h36 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_54 : _GEN_1854; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1856 = 6'h37 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_55 : _GEN_1855; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1857 = 6'h38 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_56 : _GEN_1856; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1858 = 6'h39 == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_57 : _GEN_1857; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1859 = 6'h3a == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_58 : _GEN_1858; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1860 = 6'h3b == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_59 : _GEN_1859; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1861 = 6'h3c == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_60 : _GEN_1860; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1862 = 6'h3d == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_61 : _GEN_1861; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1863 = 6'h3e == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_62 : _GEN_1862; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_51 = 6'h3f == _myTriMemVec2_19_T_1[5:0] ? myHhdoutVec_63 : _GEN_1863; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1866 = 6'h1 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1867 = 6'h2 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_2 : _GEN_1866; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1868 = 6'h3 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_3 : _GEN_1867; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1869 = 6'h4 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_4 : _GEN_1868; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1870 = 6'h5 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_5 : _GEN_1869; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1871 = 6'h6 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_6 : _GEN_1870; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1872 = 6'h7 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_7 : _GEN_1871; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1873 = 6'h8 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_8 : _GEN_1872; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1874 = 6'h9 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_9 : _GEN_1873; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1875 = 6'ha == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_10 : _GEN_1874; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1876 = 6'hb == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_11 : _GEN_1875; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1877 = 6'hc == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_12 : _GEN_1876; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1878 = 6'hd == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_13 : _GEN_1877; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1879 = 6'he == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_14 : _GEN_1878; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1880 = 6'hf == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_15 : _GEN_1879; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1881 = 6'h10 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_16 : _GEN_1880; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1882 = 6'h11 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_17 : _GEN_1881; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1883 = 6'h12 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_18 : _GEN_1882; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1884 = 6'h13 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_19 : _GEN_1883; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1885 = 6'h14 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_20 : _GEN_1884; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1886 = 6'h15 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_21 : _GEN_1885; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1887 = 6'h16 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_22 : _GEN_1886; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1888 = 6'h17 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_23 : _GEN_1887; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1889 = 6'h18 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_24 : _GEN_1888; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1890 = 6'h19 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_25 : _GEN_1889; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1891 = 6'h1a == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_26 : _GEN_1890; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1892 = 6'h1b == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_27 : _GEN_1891; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1893 = 6'h1c == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_28 : _GEN_1892; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1894 = 6'h1d == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_29 : _GEN_1893; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1895 = 6'h1e == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_30 : _GEN_1894; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1896 = 6'h1f == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_31 : _GEN_1895; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1897 = 6'h20 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_32 : _GEN_1896; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1898 = 6'h21 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_33 : _GEN_1897; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1899 = 6'h22 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_34 : _GEN_1898; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1900 = 6'h23 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_35 : _GEN_1899; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1901 = 6'h24 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_36 : _GEN_1900; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1902 = 6'h25 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_37 : _GEN_1901; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1903 = 6'h26 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_38 : _GEN_1902; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1904 = 6'h27 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_39 : _GEN_1903; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1905 = 6'h28 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_40 : _GEN_1904; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1906 = 6'h29 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_41 : _GEN_1905; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1907 = 6'h2a == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_42 : _GEN_1906; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1908 = 6'h2b == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_43 : _GEN_1907; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1909 = 6'h2c == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_44 : _GEN_1908; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1910 = 6'h2d == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_45 : _GEN_1909; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1911 = 6'h2e == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_46 : _GEN_1910; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1912 = 6'h2f == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_47 : _GEN_1911; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1913 = 6'h30 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_48 : _GEN_1912; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1914 = 6'h31 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_49 : _GEN_1913; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1915 = 6'h32 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_50 : _GEN_1914; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1916 = 6'h33 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_51 : _GEN_1915; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1917 = 6'h34 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_52 : _GEN_1916; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1918 = 6'h35 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_53 : _GEN_1917; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1919 = 6'h36 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_54 : _GEN_1918; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1920 = 6'h37 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_55 : _GEN_1919; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1921 = 6'h38 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_56 : _GEN_1920; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1922 = 6'h39 == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_57 : _GEN_1921; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1923 = 6'h3a == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_58 : _GEN_1922; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1924 = 6'h3b == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_59 : _GEN_1923; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1925 = 6'h3c == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_60 : _GEN_1924; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1926 = 6'h3d == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_61 : _GEN_1925; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1927 = 6'h3e == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_62 : _GEN_1926; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_50 = 6'h3f == _myTriMemVec2_18_T_1[5:0] ? myHhdoutVec_63 : _GEN_1927; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1930 = 6'h1 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1931 = 6'h2 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_2 : _GEN_1930; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1932 = 6'h3 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_3 : _GEN_1931; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1933 = 6'h4 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_4 : _GEN_1932; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1934 = 6'h5 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_5 : _GEN_1933; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1935 = 6'h6 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_6 : _GEN_1934; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1936 = 6'h7 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_7 : _GEN_1935; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1937 = 6'h8 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_8 : _GEN_1936; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1938 = 6'h9 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_9 : _GEN_1937; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1939 = 6'ha == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_10 : _GEN_1938; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1940 = 6'hb == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_11 : _GEN_1939; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1941 = 6'hc == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_12 : _GEN_1940; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1942 = 6'hd == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_13 : _GEN_1941; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1943 = 6'he == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_14 : _GEN_1942; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1944 = 6'hf == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_15 : _GEN_1943; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1945 = 6'h10 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_16 : _GEN_1944; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1946 = 6'h11 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_17 : _GEN_1945; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1947 = 6'h12 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_18 : _GEN_1946; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1948 = 6'h13 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_19 : _GEN_1947; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1949 = 6'h14 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_20 : _GEN_1948; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1950 = 6'h15 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_21 : _GEN_1949; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1951 = 6'h16 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_22 : _GEN_1950; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1952 = 6'h17 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_23 : _GEN_1951; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1953 = 6'h18 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_24 : _GEN_1952; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1954 = 6'h19 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_25 : _GEN_1953; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1955 = 6'h1a == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_26 : _GEN_1954; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1956 = 6'h1b == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_27 : _GEN_1955; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1957 = 6'h1c == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_28 : _GEN_1956; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1958 = 6'h1d == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_29 : _GEN_1957; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1959 = 6'h1e == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_30 : _GEN_1958; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1960 = 6'h1f == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_31 : _GEN_1959; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1961 = 6'h20 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_32 : _GEN_1960; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1962 = 6'h21 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_33 : _GEN_1961; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1963 = 6'h22 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_34 : _GEN_1962; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1964 = 6'h23 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_35 : _GEN_1963; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1965 = 6'h24 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_36 : _GEN_1964; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1966 = 6'h25 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_37 : _GEN_1965; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1967 = 6'h26 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_38 : _GEN_1966; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1968 = 6'h27 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_39 : _GEN_1967; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1969 = 6'h28 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_40 : _GEN_1968; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1970 = 6'h29 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_41 : _GEN_1969; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1971 = 6'h2a == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_42 : _GEN_1970; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1972 = 6'h2b == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_43 : _GEN_1971; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1973 = 6'h2c == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_44 : _GEN_1972; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1974 = 6'h2d == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_45 : _GEN_1973; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1975 = 6'h2e == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_46 : _GEN_1974; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1976 = 6'h2f == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_47 : _GEN_1975; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1977 = 6'h30 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_48 : _GEN_1976; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1978 = 6'h31 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_49 : _GEN_1977; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1979 = 6'h32 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_50 : _GEN_1978; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1980 = 6'h33 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_51 : _GEN_1979; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1981 = 6'h34 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_52 : _GEN_1980; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1982 = 6'h35 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_53 : _GEN_1981; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1983 = 6'h36 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_54 : _GEN_1982; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1984 = 6'h37 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_55 : _GEN_1983; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1985 = 6'h38 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_56 : _GEN_1984; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1986 = 6'h39 == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_57 : _GEN_1985; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1987 = 6'h3a == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_58 : _GEN_1986; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1988 = 6'h3b == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_59 : _GEN_1987; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1989 = 6'h3c == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_60 : _GEN_1988; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1990 = 6'h3d == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_61 : _GEN_1989; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1991 = 6'h3e == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_62 : _GEN_1990; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_49 = 6'h3f == _myTriMemVec2_17_T_1[5:0] ? myHhdoutVec_63 : _GEN_1991; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1994 = 6'h1 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1995 = 6'h2 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_2 : _GEN_1994; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1996 = 6'h3 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_3 : _GEN_1995; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1997 = 6'h4 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_4 : _GEN_1996; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1998 = 6'h5 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_5 : _GEN_1997; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_1999 = 6'h6 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_6 : _GEN_1998; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2000 = 6'h7 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_7 : _GEN_1999; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2001 = 6'h8 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_8 : _GEN_2000; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2002 = 6'h9 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_9 : _GEN_2001; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2003 = 6'ha == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_10 : _GEN_2002; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2004 = 6'hb == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_11 : _GEN_2003; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2005 = 6'hc == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_12 : _GEN_2004; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2006 = 6'hd == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_13 : _GEN_2005; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2007 = 6'he == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_14 : _GEN_2006; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2008 = 6'hf == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_15 : _GEN_2007; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2009 = 6'h10 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_16 : _GEN_2008; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2010 = 6'h11 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_17 : _GEN_2009; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2011 = 6'h12 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_18 : _GEN_2010; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2012 = 6'h13 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_19 : _GEN_2011; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2013 = 6'h14 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_20 : _GEN_2012; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2014 = 6'h15 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_21 : _GEN_2013; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2015 = 6'h16 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_22 : _GEN_2014; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2016 = 6'h17 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_23 : _GEN_2015; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2017 = 6'h18 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_24 : _GEN_2016; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2018 = 6'h19 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_25 : _GEN_2017; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2019 = 6'h1a == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_26 : _GEN_2018; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2020 = 6'h1b == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_27 : _GEN_2019; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2021 = 6'h1c == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_28 : _GEN_2020; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2022 = 6'h1d == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_29 : _GEN_2021; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2023 = 6'h1e == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_30 : _GEN_2022; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2024 = 6'h1f == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_31 : _GEN_2023; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2025 = 6'h20 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_32 : _GEN_2024; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2026 = 6'h21 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_33 : _GEN_2025; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2027 = 6'h22 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_34 : _GEN_2026; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2028 = 6'h23 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_35 : _GEN_2027; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2029 = 6'h24 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_36 : _GEN_2028; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2030 = 6'h25 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_37 : _GEN_2029; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2031 = 6'h26 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_38 : _GEN_2030; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2032 = 6'h27 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_39 : _GEN_2031; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2033 = 6'h28 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_40 : _GEN_2032; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2034 = 6'h29 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_41 : _GEN_2033; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2035 = 6'h2a == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_42 : _GEN_2034; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2036 = 6'h2b == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_43 : _GEN_2035; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2037 = 6'h2c == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_44 : _GEN_2036; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2038 = 6'h2d == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_45 : _GEN_2037; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2039 = 6'h2e == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_46 : _GEN_2038; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2040 = 6'h2f == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_47 : _GEN_2039; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2041 = 6'h30 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_48 : _GEN_2040; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2042 = 6'h31 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_49 : _GEN_2041; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2043 = 6'h32 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_50 : _GEN_2042; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2044 = 6'h33 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_51 : _GEN_2043; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2045 = 6'h34 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_52 : _GEN_2044; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2046 = 6'h35 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_53 : _GEN_2045; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2047 = 6'h36 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_54 : _GEN_2046; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2048 = 6'h37 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_55 : _GEN_2047; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2049 = 6'h38 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_56 : _GEN_2048; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2050 = 6'h39 == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_57 : _GEN_2049; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2051 = 6'h3a == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_58 : _GEN_2050; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2052 = 6'h3b == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_59 : _GEN_2051; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2053 = 6'h3c == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_60 : _GEN_2052; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2054 = 6'h3d == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_61 : _GEN_2053; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2055 = 6'h3e == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_62 : _GEN_2054; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_48 = 6'h3f == _myTriMemVec2_16_T_1[5:0] ? myHhdoutVec_63 : _GEN_2055; // @[hh_core.scala 149:{52,52}]
  wire [255:0] myHhdoutWire_hi_hi_lo = {myHhdoutVec2_55,myHhdoutVec2_54,myHhdoutVec2_53,myHhdoutVec2_52,myHhdoutVec2_51,
    myHhdoutVec2_50,myHhdoutVec2_49,myHhdoutVec2_48}; // @[hh_core.scala 153:42]
  wire [31:0] _GEN_2058 = 6'h1 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2059 = 6'h2 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_2 : _GEN_2058; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2060 = 6'h3 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_3 : _GEN_2059; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2061 = 6'h4 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_4 : _GEN_2060; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2062 = 6'h5 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_5 : _GEN_2061; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2063 = 6'h6 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_6 : _GEN_2062; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2064 = 6'h7 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_7 : _GEN_2063; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2065 = 6'h8 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_8 : _GEN_2064; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2066 = 6'h9 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_9 : _GEN_2065; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2067 = 6'ha == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_10 : _GEN_2066; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2068 = 6'hb == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_11 : _GEN_2067; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2069 = 6'hc == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_12 : _GEN_2068; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2070 = 6'hd == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_13 : _GEN_2069; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2071 = 6'he == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_14 : _GEN_2070; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2072 = 6'hf == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_15 : _GEN_2071; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2073 = 6'h10 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_16 : _GEN_2072; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2074 = 6'h11 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_17 : _GEN_2073; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2075 = 6'h12 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_18 : _GEN_2074; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2076 = 6'h13 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_19 : _GEN_2075; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2077 = 6'h14 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_20 : _GEN_2076; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2078 = 6'h15 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_21 : _GEN_2077; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2079 = 6'h16 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_22 : _GEN_2078; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2080 = 6'h17 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_23 : _GEN_2079; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2081 = 6'h18 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_24 : _GEN_2080; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2082 = 6'h19 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_25 : _GEN_2081; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2083 = 6'h1a == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_26 : _GEN_2082; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2084 = 6'h1b == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_27 : _GEN_2083; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2085 = 6'h1c == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_28 : _GEN_2084; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2086 = 6'h1d == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_29 : _GEN_2085; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2087 = 6'h1e == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_30 : _GEN_2086; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2088 = 6'h1f == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_31 : _GEN_2087; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2089 = 6'h20 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_32 : _GEN_2088; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2090 = 6'h21 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_33 : _GEN_2089; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2091 = 6'h22 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_34 : _GEN_2090; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2092 = 6'h23 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_35 : _GEN_2091; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2093 = 6'h24 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_36 : _GEN_2092; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2094 = 6'h25 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_37 : _GEN_2093; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2095 = 6'h26 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_38 : _GEN_2094; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2096 = 6'h27 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_39 : _GEN_2095; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2097 = 6'h28 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_40 : _GEN_2096; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2098 = 6'h29 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_41 : _GEN_2097; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2099 = 6'h2a == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_42 : _GEN_2098; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2100 = 6'h2b == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_43 : _GEN_2099; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2101 = 6'h2c == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_44 : _GEN_2100; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2102 = 6'h2d == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_45 : _GEN_2101; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2103 = 6'h2e == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_46 : _GEN_2102; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2104 = 6'h2f == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_47 : _GEN_2103; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2105 = 6'h30 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_48 : _GEN_2104; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2106 = 6'h31 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_49 : _GEN_2105; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2107 = 6'h32 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_50 : _GEN_2106; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2108 = 6'h33 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_51 : _GEN_2107; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2109 = 6'h34 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_52 : _GEN_2108; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2110 = 6'h35 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_53 : _GEN_2109; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2111 = 6'h36 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_54 : _GEN_2110; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2112 = 6'h37 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_55 : _GEN_2111; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2113 = 6'h38 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_56 : _GEN_2112; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2114 = 6'h39 == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_57 : _GEN_2113; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2115 = 6'h3a == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_58 : _GEN_2114; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2116 = 6'h3b == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_59 : _GEN_2115; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2117 = 6'h3c == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_60 : _GEN_2116; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2118 = 6'h3d == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_61 : _GEN_2117; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2119 = 6'h3e == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_62 : _GEN_2118; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_47 = 6'h3f == _myTriMemVec2_15_T_1[5:0] ? myHhdoutVec_63 : _GEN_2119; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2122 = 6'h1 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2123 = 6'h2 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_2 : _GEN_2122; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2124 = 6'h3 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_3 : _GEN_2123; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2125 = 6'h4 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_4 : _GEN_2124; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2126 = 6'h5 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_5 : _GEN_2125; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2127 = 6'h6 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_6 : _GEN_2126; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2128 = 6'h7 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_7 : _GEN_2127; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2129 = 6'h8 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_8 : _GEN_2128; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2130 = 6'h9 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_9 : _GEN_2129; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2131 = 6'ha == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_10 : _GEN_2130; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2132 = 6'hb == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_11 : _GEN_2131; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2133 = 6'hc == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_12 : _GEN_2132; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2134 = 6'hd == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_13 : _GEN_2133; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2135 = 6'he == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_14 : _GEN_2134; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2136 = 6'hf == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_15 : _GEN_2135; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2137 = 6'h10 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_16 : _GEN_2136; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2138 = 6'h11 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_17 : _GEN_2137; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2139 = 6'h12 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_18 : _GEN_2138; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2140 = 6'h13 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_19 : _GEN_2139; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2141 = 6'h14 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_20 : _GEN_2140; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2142 = 6'h15 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_21 : _GEN_2141; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2143 = 6'h16 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_22 : _GEN_2142; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2144 = 6'h17 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_23 : _GEN_2143; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2145 = 6'h18 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_24 : _GEN_2144; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2146 = 6'h19 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_25 : _GEN_2145; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2147 = 6'h1a == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_26 : _GEN_2146; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2148 = 6'h1b == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_27 : _GEN_2147; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2149 = 6'h1c == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_28 : _GEN_2148; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2150 = 6'h1d == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_29 : _GEN_2149; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2151 = 6'h1e == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_30 : _GEN_2150; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2152 = 6'h1f == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_31 : _GEN_2151; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2153 = 6'h20 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_32 : _GEN_2152; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2154 = 6'h21 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_33 : _GEN_2153; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2155 = 6'h22 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_34 : _GEN_2154; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2156 = 6'h23 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_35 : _GEN_2155; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2157 = 6'h24 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_36 : _GEN_2156; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2158 = 6'h25 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_37 : _GEN_2157; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2159 = 6'h26 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_38 : _GEN_2158; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2160 = 6'h27 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_39 : _GEN_2159; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2161 = 6'h28 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_40 : _GEN_2160; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2162 = 6'h29 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_41 : _GEN_2161; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2163 = 6'h2a == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_42 : _GEN_2162; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2164 = 6'h2b == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_43 : _GEN_2163; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2165 = 6'h2c == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_44 : _GEN_2164; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2166 = 6'h2d == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_45 : _GEN_2165; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2167 = 6'h2e == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_46 : _GEN_2166; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2168 = 6'h2f == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_47 : _GEN_2167; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2169 = 6'h30 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_48 : _GEN_2168; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2170 = 6'h31 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_49 : _GEN_2169; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2171 = 6'h32 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_50 : _GEN_2170; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2172 = 6'h33 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_51 : _GEN_2171; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2173 = 6'h34 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_52 : _GEN_2172; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2174 = 6'h35 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_53 : _GEN_2173; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2175 = 6'h36 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_54 : _GEN_2174; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2176 = 6'h37 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_55 : _GEN_2175; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2177 = 6'h38 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_56 : _GEN_2176; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2178 = 6'h39 == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_57 : _GEN_2177; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2179 = 6'h3a == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_58 : _GEN_2178; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2180 = 6'h3b == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_59 : _GEN_2179; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2181 = 6'h3c == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_60 : _GEN_2180; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2182 = 6'h3d == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_61 : _GEN_2181; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2183 = 6'h3e == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_62 : _GEN_2182; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_46 = 6'h3f == _myTriMemVec2_14_T_1[5:0] ? myHhdoutVec_63 : _GEN_2183; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2186 = 6'h1 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2187 = 6'h2 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_2 : _GEN_2186; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2188 = 6'h3 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_3 : _GEN_2187; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2189 = 6'h4 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_4 : _GEN_2188; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2190 = 6'h5 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_5 : _GEN_2189; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2191 = 6'h6 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_6 : _GEN_2190; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2192 = 6'h7 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_7 : _GEN_2191; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2193 = 6'h8 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_8 : _GEN_2192; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2194 = 6'h9 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_9 : _GEN_2193; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2195 = 6'ha == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_10 : _GEN_2194; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2196 = 6'hb == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_11 : _GEN_2195; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2197 = 6'hc == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_12 : _GEN_2196; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2198 = 6'hd == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_13 : _GEN_2197; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2199 = 6'he == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_14 : _GEN_2198; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2200 = 6'hf == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_15 : _GEN_2199; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2201 = 6'h10 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_16 : _GEN_2200; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2202 = 6'h11 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_17 : _GEN_2201; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2203 = 6'h12 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_18 : _GEN_2202; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2204 = 6'h13 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_19 : _GEN_2203; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2205 = 6'h14 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_20 : _GEN_2204; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2206 = 6'h15 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_21 : _GEN_2205; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2207 = 6'h16 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_22 : _GEN_2206; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2208 = 6'h17 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_23 : _GEN_2207; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2209 = 6'h18 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_24 : _GEN_2208; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2210 = 6'h19 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_25 : _GEN_2209; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2211 = 6'h1a == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_26 : _GEN_2210; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2212 = 6'h1b == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_27 : _GEN_2211; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2213 = 6'h1c == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_28 : _GEN_2212; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2214 = 6'h1d == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_29 : _GEN_2213; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2215 = 6'h1e == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_30 : _GEN_2214; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2216 = 6'h1f == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_31 : _GEN_2215; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2217 = 6'h20 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_32 : _GEN_2216; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2218 = 6'h21 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_33 : _GEN_2217; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2219 = 6'h22 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_34 : _GEN_2218; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2220 = 6'h23 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_35 : _GEN_2219; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2221 = 6'h24 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_36 : _GEN_2220; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2222 = 6'h25 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_37 : _GEN_2221; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2223 = 6'h26 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_38 : _GEN_2222; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2224 = 6'h27 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_39 : _GEN_2223; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2225 = 6'h28 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_40 : _GEN_2224; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2226 = 6'h29 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_41 : _GEN_2225; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2227 = 6'h2a == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_42 : _GEN_2226; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2228 = 6'h2b == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_43 : _GEN_2227; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2229 = 6'h2c == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_44 : _GEN_2228; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2230 = 6'h2d == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_45 : _GEN_2229; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2231 = 6'h2e == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_46 : _GEN_2230; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2232 = 6'h2f == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_47 : _GEN_2231; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2233 = 6'h30 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_48 : _GEN_2232; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2234 = 6'h31 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_49 : _GEN_2233; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2235 = 6'h32 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_50 : _GEN_2234; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2236 = 6'h33 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_51 : _GEN_2235; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2237 = 6'h34 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_52 : _GEN_2236; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2238 = 6'h35 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_53 : _GEN_2237; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2239 = 6'h36 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_54 : _GEN_2238; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2240 = 6'h37 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_55 : _GEN_2239; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2241 = 6'h38 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_56 : _GEN_2240; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2242 = 6'h39 == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_57 : _GEN_2241; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2243 = 6'h3a == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_58 : _GEN_2242; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2244 = 6'h3b == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_59 : _GEN_2243; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2245 = 6'h3c == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_60 : _GEN_2244; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2246 = 6'h3d == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_61 : _GEN_2245; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2247 = 6'h3e == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_62 : _GEN_2246; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_45 = 6'h3f == _myTriMemVec2_13_T_1[5:0] ? myHhdoutVec_63 : _GEN_2247; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2250 = 6'h1 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2251 = 6'h2 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_2 : _GEN_2250; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2252 = 6'h3 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_3 : _GEN_2251; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2253 = 6'h4 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_4 : _GEN_2252; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2254 = 6'h5 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_5 : _GEN_2253; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2255 = 6'h6 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_6 : _GEN_2254; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2256 = 6'h7 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_7 : _GEN_2255; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2257 = 6'h8 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_8 : _GEN_2256; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2258 = 6'h9 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_9 : _GEN_2257; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2259 = 6'ha == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_10 : _GEN_2258; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2260 = 6'hb == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_11 : _GEN_2259; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2261 = 6'hc == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_12 : _GEN_2260; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2262 = 6'hd == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_13 : _GEN_2261; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2263 = 6'he == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_14 : _GEN_2262; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2264 = 6'hf == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_15 : _GEN_2263; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2265 = 6'h10 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_16 : _GEN_2264; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2266 = 6'h11 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_17 : _GEN_2265; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2267 = 6'h12 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_18 : _GEN_2266; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2268 = 6'h13 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_19 : _GEN_2267; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2269 = 6'h14 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_20 : _GEN_2268; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2270 = 6'h15 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_21 : _GEN_2269; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2271 = 6'h16 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_22 : _GEN_2270; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2272 = 6'h17 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_23 : _GEN_2271; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2273 = 6'h18 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_24 : _GEN_2272; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2274 = 6'h19 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_25 : _GEN_2273; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2275 = 6'h1a == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_26 : _GEN_2274; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2276 = 6'h1b == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_27 : _GEN_2275; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2277 = 6'h1c == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_28 : _GEN_2276; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2278 = 6'h1d == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_29 : _GEN_2277; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2279 = 6'h1e == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_30 : _GEN_2278; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2280 = 6'h1f == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_31 : _GEN_2279; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2281 = 6'h20 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_32 : _GEN_2280; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2282 = 6'h21 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_33 : _GEN_2281; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2283 = 6'h22 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_34 : _GEN_2282; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2284 = 6'h23 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_35 : _GEN_2283; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2285 = 6'h24 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_36 : _GEN_2284; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2286 = 6'h25 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_37 : _GEN_2285; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2287 = 6'h26 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_38 : _GEN_2286; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2288 = 6'h27 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_39 : _GEN_2287; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2289 = 6'h28 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_40 : _GEN_2288; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2290 = 6'h29 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_41 : _GEN_2289; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2291 = 6'h2a == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_42 : _GEN_2290; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2292 = 6'h2b == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_43 : _GEN_2291; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2293 = 6'h2c == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_44 : _GEN_2292; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2294 = 6'h2d == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_45 : _GEN_2293; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2295 = 6'h2e == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_46 : _GEN_2294; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2296 = 6'h2f == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_47 : _GEN_2295; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2297 = 6'h30 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_48 : _GEN_2296; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2298 = 6'h31 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_49 : _GEN_2297; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2299 = 6'h32 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_50 : _GEN_2298; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2300 = 6'h33 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_51 : _GEN_2299; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2301 = 6'h34 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_52 : _GEN_2300; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2302 = 6'h35 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_53 : _GEN_2301; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2303 = 6'h36 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_54 : _GEN_2302; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2304 = 6'h37 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_55 : _GEN_2303; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2305 = 6'h38 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_56 : _GEN_2304; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2306 = 6'h39 == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_57 : _GEN_2305; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2307 = 6'h3a == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_58 : _GEN_2306; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2308 = 6'h3b == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_59 : _GEN_2307; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2309 = 6'h3c == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_60 : _GEN_2308; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2310 = 6'h3d == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_61 : _GEN_2309; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2311 = 6'h3e == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_62 : _GEN_2310; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_44 = 6'h3f == _myTriMemVec2_12_T_1[5:0] ? myHhdoutVec_63 : _GEN_2311; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2314 = 6'h1 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2315 = 6'h2 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_2 : _GEN_2314; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2316 = 6'h3 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_3 : _GEN_2315; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2317 = 6'h4 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_4 : _GEN_2316; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2318 = 6'h5 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_5 : _GEN_2317; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2319 = 6'h6 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_6 : _GEN_2318; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2320 = 6'h7 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_7 : _GEN_2319; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2321 = 6'h8 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_8 : _GEN_2320; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2322 = 6'h9 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_9 : _GEN_2321; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2323 = 6'ha == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_10 : _GEN_2322; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2324 = 6'hb == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_11 : _GEN_2323; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2325 = 6'hc == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_12 : _GEN_2324; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2326 = 6'hd == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_13 : _GEN_2325; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2327 = 6'he == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_14 : _GEN_2326; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2328 = 6'hf == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_15 : _GEN_2327; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2329 = 6'h10 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_16 : _GEN_2328; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2330 = 6'h11 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_17 : _GEN_2329; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2331 = 6'h12 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_18 : _GEN_2330; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2332 = 6'h13 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_19 : _GEN_2331; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2333 = 6'h14 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_20 : _GEN_2332; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2334 = 6'h15 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_21 : _GEN_2333; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2335 = 6'h16 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_22 : _GEN_2334; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2336 = 6'h17 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_23 : _GEN_2335; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2337 = 6'h18 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_24 : _GEN_2336; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2338 = 6'h19 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_25 : _GEN_2337; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2339 = 6'h1a == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_26 : _GEN_2338; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2340 = 6'h1b == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_27 : _GEN_2339; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2341 = 6'h1c == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_28 : _GEN_2340; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2342 = 6'h1d == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_29 : _GEN_2341; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2343 = 6'h1e == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_30 : _GEN_2342; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2344 = 6'h1f == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_31 : _GEN_2343; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2345 = 6'h20 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_32 : _GEN_2344; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2346 = 6'h21 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_33 : _GEN_2345; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2347 = 6'h22 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_34 : _GEN_2346; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2348 = 6'h23 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_35 : _GEN_2347; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2349 = 6'h24 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_36 : _GEN_2348; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2350 = 6'h25 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_37 : _GEN_2349; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2351 = 6'h26 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_38 : _GEN_2350; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2352 = 6'h27 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_39 : _GEN_2351; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2353 = 6'h28 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_40 : _GEN_2352; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2354 = 6'h29 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_41 : _GEN_2353; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2355 = 6'h2a == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_42 : _GEN_2354; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2356 = 6'h2b == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_43 : _GEN_2355; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2357 = 6'h2c == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_44 : _GEN_2356; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2358 = 6'h2d == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_45 : _GEN_2357; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2359 = 6'h2e == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_46 : _GEN_2358; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2360 = 6'h2f == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_47 : _GEN_2359; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2361 = 6'h30 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_48 : _GEN_2360; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2362 = 6'h31 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_49 : _GEN_2361; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2363 = 6'h32 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_50 : _GEN_2362; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2364 = 6'h33 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_51 : _GEN_2363; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2365 = 6'h34 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_52 : _GEN_2364; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2366 = 6'h35 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_53 : _GEN_2365; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2367 = 6'h36 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_54 : _GEN_2366; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2368 = 6'h37 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_55 : _GEN_2367; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2369 = 6'h38 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_56 : _GEN_2368; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2370 = 6'h39 == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_57 : _GEN_2369; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2371 = 6'h3a == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_58 : _GEN_2370; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2372 = 6'h3b == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_59 : _GEN_2371; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2373 = 6'h3c == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_60 : _GEN_2372; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2374 = 6'h3d == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_61 : _GEN_2373; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2375 = 6'h3e == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_62 : _GEN_2374; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_43 = 6'h3f == _myTriMemVec2_11_T_1[5:0] ? myHhdoutVec_63 : _GEN_2375; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2378 = 6'h1 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2379 = 6'h2 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_2 : _GEN_2378; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2380 = 6'h3 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_3 : _GEN_2379; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2381 = 6'h4 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_4 : _GEN_2380; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2382 = 6'h5 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_5 : _GEN_2381; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2383 = 6'h6 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_6 : _GEN_2382; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2384 = 6'h7 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_7 : _GEN_2383; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2385 = 6'h8 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_8 : _GEN_2384; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2386 = 6'h9 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_9 : _GEN_2385; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2387 = 6'ha == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_10 : _GEN_2386; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2388 = 6'hb == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_11 : _GEN_2387; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2389 = 6'hc == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_12 : _GEN_2388; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2390 = 6'hd == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_13 : _GEN_2389; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2391 = 6'he == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_14 : _GEN_2390; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2392 = 6'hf == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_15 : _GEN_2391; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2393 = 6'h10 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_16 : _GEN_2392; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2394 = 6'h11 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_17 : _GEN_2393; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2395 = 6'h12 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_18 : _GEN_2394; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2396 = 6'h13 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_19 : _GEN_2395; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2397 = 6'h14 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_20 : _GEN_2396; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2398 = 6'h15 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_21 : _GEN_2397; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2399 = 6'h16 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_22 : _GEN_2398; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2400 = 6'h17 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_23 : _GEN_2399; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2401 = 6'h18 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_24 : _GEN_2400; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2402 = 6'h19 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_25 : _GEN_2401; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2403 = 6'h1a == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_26 : _GEN_2402; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2404 = 6'h1b == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_27 : _GEN_2403; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2405 = 6'h1c == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_28 : _GEN_2404; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2406 = 6'h1d == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_29 : _GEN_2405; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2407 = 6'h1e == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_30 : _GEN_2406; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2408 = 6'h1f == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_31 : _GEN_2407; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2409 = 6'h20 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_32 : _GEN_2408; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2410 = 6'h21 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_33 : _GEN_2409; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2411 = 6'h22 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_34 : _GEN_2410; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2412 = 6'h23 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_35 : _GEN_2411; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2413 = 6'h24 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_36 : _GEN_2412; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2414 = 6'h25 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_37 : _GEN_2413; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2415 = 6'h26 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_38 : _GEN_2414; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2416 = 6'h27 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_39 : _GEN_2415; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2417 = 6'h28 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_40 : _GEN_2416; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2418 = 6'h29 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_41 : _GEN_2417; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2419 = 6'h2a == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_42 : _GEN_2418; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2420 = 6'h2b == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_43 : _GEN_2419; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2421 = 6'h2c == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_44 : _GEN_2420; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2422 = 6'h2d == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_45 : _GEN_2421; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2423 = 6'h2e == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_46 : _GEN_2422; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2424 = 6'h2f == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_47 : _GEN_2423; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2425 = 6'h30 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_48 : _GEN_2424; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2426 = 6'h31 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_49 : _GEN_2425; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2427 = 6'h32 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_50 : _GEN_2426; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2428 = 6'h33 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_51 : _GEN_2427; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2429 = 6'h34 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_52 : _GEN_2428; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2430 = 6'h35 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_53 : _GEN_2429; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2431 = 6'h36 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_54 : _GEN_2430; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2432 = 6'h37 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_55 : _GEN_2431; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2433 = 6'h38 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_56 : _GEN_2432; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2434 = 6'h39 == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_57 : _GEN_2433; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2435 = 6'h3a == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_58 : _GEN_2434; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2436 = 6'h3b == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_59 : _GEN_2435; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2437 = 6'h3c == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_60 : _GEN_2436; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2438 = 6'h3d == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_61 : _GEN_2437; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2439 = 6'h3e == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_62 : _GEN_2438; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_42 = 6'h3f == _myTriMemVec2_10_T_1[5:0] ? myHhdoutVec_63 : _GEN_2439; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2442 = 6'h1 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2443 = 6'h2 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_2 : _GEN_2442; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2444 = 6'h3 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_3 : _GEN_2443; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2445 = 6'h4 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_4 : _GEN_2444; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2446 = 6'h5 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_5 : _GEN_2445; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2447 = 6'h6 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_6 : _GEN_2446; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2448 = 6'h7 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_7 : _GEN_2447; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2449 = 6'h8 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_8 : _GEN_2448; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2450 = 6'h9 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_9 : _GEN_2449; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2451 = 6'ha == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_10 : _GEN_2450; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2452 = 6'hb == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_11 : _GEN_2451; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2453 = 6'hc == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_12 : _GEN_2452; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2454 = 6'hd == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_13 : _GEN_2453; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2455 = 6'he == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_14 : _GEN_2454; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2456 = 6'hf == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_15 : _GEN_2455; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2457 = 6'h10 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_16 : _GEN_2456; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2458 = 6'h11 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_17 : _GEN_2457; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2459 = 6'h12 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_18 : _GEN_2458; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2460 = 6'h13 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_19 : _GEN_2459; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2461 = 6'h14 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_20 : _GEN_2460; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2462 = 6'h15 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_21 : _GEN_2461; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2463 = 6'h16 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_22 : _GEN_2462; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2464 = 6'h17 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_23 : _GEN_2463; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2465 = 6'h18 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_24 : _GEN_2464; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2466 = 6'h19 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_25 : _GEN_2465; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2467 = 6'h1a == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_26 : _GEN_2466; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2468 = 6'h1b == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_27 : _GEN_2467; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2469 = 6'h1c == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_28 : _GEN_2468; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2470 = 6'h1d == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_29 : _GEN_2469; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2471 = 6'h1e == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_30 : _GEN_2470; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2472 = 6'h1f == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_31 : _GEN_2471; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2473 = 6'h20 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_32 : _GEN_2472; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2474 = 6'h21 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_33 : _GEN_2473; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2475 = 6'h22 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_34 : _GEN_2474; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2476 = 6'h23 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_35 : _GEN_2475; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2477 = 6'h24 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_36 : _GEN_2476; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2478 = 6'h25 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_37 : _GEN_2477; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2479 = 6'h26 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_38 : _GEN_2478; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2480 = 6'h27 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_39 : _GEN_2479; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2481 = 6'h28 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_40 : _GEN_2480; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2482 = 6'h29 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_41 : _GEN_2481; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2483 = 6'h2a == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_42 : _GEN_2482; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2484 = 6'h2b == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_43 : _GEN_2483; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2485 = 6'h2c == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_44 : _GEN_2484; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2486 = 6'h2d == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_45 : _GEN_2485; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2487 = 6'h2e == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_46 : _GEN_2486; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2488 = 6'h2f == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_47 : _GEN_2487; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2489 = 6'h30 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_48 : _GEN_2488; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2490 = 6'h31 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_49 : _GEN_2489; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2491 = 6'h32 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_50 : _GEN_2490; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2492 = 6'h33 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_51 : _GEN_2491; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2493 = 6'h34 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_52 : _GEN_2492; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2494 = 6'h35 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_53 : _GEN_2493; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2495 = 6'h36 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_54 : _GEN_2494; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2496 = 6'h37 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_55 : _GEN_2495; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2497 = 6'h38 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_56 : _GEN_2496; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2498 = 6'h39 == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_57 : _GEN_2497; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2499 = 6'h3a == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_58 : _GEN_2498; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2500 = 6'h3b == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_59 : _GEN_2499; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2501 = 6'h3c == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_60 : _GEN_2500; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2502 = 6'h3d == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_61 : _GEN_2501; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2503 = 6'h3e == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_62 : _GEN_2502; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_41 = 6'h3f == _myTriMemVec2_9_T_1[5:0] ? myHhdoutVec_63 : _GEN_2503; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2506 = 6'h1 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2507 = 6'h2 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_2 : _GEN_2506; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2508 = 6'h3 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_3 : _GEN_2507; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2509 = 6'h4 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_4 : _GEN_2508; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2510 = 6'h5 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_5 : _GEN_2509; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2511 = 6'h6 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_6 : _GEN_2510; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2512 = 6'h7 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_7 : _GEN_2511; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2513 = 6'h8 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_8 : _GEN_2512; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2514 = 6'h9 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_9 : _GEN_2513; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2515 = 6'ha == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_10 : _GEN_2514; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2516 = 6'hb == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_11 : _GEN_2515; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2517 = 6'hc == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_12 : _GEN_2516; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2518 = 6'hd == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_13 : _GEN_2517; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2519 = 6'he == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_14 : _GEN_2518; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2520 = 6'hf == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_15 : _GEN_2519; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2521 = 6'h10 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_16 : _GEN_2520; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2522 = 6'h11 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_17 : _GEN_2521; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2523 = 6'h12 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_18 : _GEN_2522; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2524 = 6'h13 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_19 : _GEN_2523; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2525 = 6'h14 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_20 : _GEN_2524; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2526 = 6'h15 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_21 : _GEN_2525; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2527 = 6'h16 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_22 : _GEN_2526; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2528 = 6'h17 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_23 : _GEN_2527; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2529 = 6'h18 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_24 : _GEN_2528; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2530 = 6'h19 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_25 : _GEN_2529; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2531 = 6'h1a == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_26 : _GEN_2530; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2532 = 6'h1b == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_27 : _GEN_2531; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2533 = 6'h1c == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_28 : _GEN_2532; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2534 = 6'h1d == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_29 : _GEN_2533; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2535 = 6'h1e == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_30 : _GEN_2534; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2536 = 6'h1f == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_31 : _GEN_2535; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2537 = 6'h20 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_32 : _GEN_2536; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2538 = 6'h21 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_33 : _GEN_2537; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2539 = 6'h22 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_34 : _GEN_2538; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2540 = 6'h23 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_35 : _GEN_2539; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2541 = 6'h24 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_36 : _GEN_2540; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2542 = 6'h25 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_37 : _GEN_2541; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2543 = 6'h26 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_38 : _GEN_2542; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2544 = 6'h27 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_39 : _GEN_2543; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2545 = 6'h28 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_40 : _GEN_2544; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2546 = 6'h29 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_41 : _GEN_2545; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2547 = 6'h2a == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_42 : _GEN_2546; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2548 = 6'h2b == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_43 : _GEN_2547; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2549 = 6'h2c == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_44 : _GEN_2548; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2550 = 6'h2d == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_45 : _GEN_2549; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2551 = 6'h2e == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_46 : _GEN_2550; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2552 = 6'h2f == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_47 : _GEN_2551; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2553 = 6'h30 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_48 : _GEN_2552; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2554 = 6'h31 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_49 : _GEN_2553; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2555 = 6'h32 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_50 : _GEN_2554; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2556 = 6'h33 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_51 : _GEN_2555; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2557 = 6'h34 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_52 : _GEN_2556; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2558 = 6'h35 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_53 : _GEN_2557; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2559 = 6'h36 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_54 : _GEN_2558; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2560 = 6'h37 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_55 : _GEN_2559; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2561 = 6'h38 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_56 : _GEN_2560; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2562 = 6'h39 == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_57 : _GEN_2561; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2563 = 6'h3a == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_58 : _GEN_2562; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2564 = 6'h3b == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_59 : _GEN_2563; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2565 = 6'h3c == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_60 : _GEN_2564; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2566 = 6'h3d == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_61 : _GEN_2565; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2567 = 6'h3e == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_62 : _GEN_2566; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_40 = 6'h3f == _myTriMemVec2_8_T_1[5:0] ? myHhdoutVec_63 : _GEN_2567; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2570 = 6'h1 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2571 = 6'h2 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_2 : _GEN_2570; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2572 = 6'h3 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_3 : _GEN_2571; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2573 = 6'h4 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_4 : _GEN_2572; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2574 = 6'h5 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_5 : _GEN_2573; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2575 = 6'h6 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_6 : _GEN_2574; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2576 = 6'h7 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_7 : _GEN_2575; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2577 = 6'h8 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_8 : _GEN_2576; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2578 = 6'h9 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_9 : _GEN_2577; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2579 = 6'ha == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_10 : _GEN_2578; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2580 = 6'hb == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_11 : _GEN_2579; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2581 = 6'hc == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_12 : _GEN_2580; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2582 = 6'hd == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_13 : _GEN_2581; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2583 = 6'he == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_14 : _GEN_2582; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2584 = 6'hf == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_15 : _GEN_2583; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2585 = 6'h10 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_16 : _GEN_2584; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2586 = 6'h11 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_17 : _GEN_2585; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2587 = 6'h12 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_18 : _GEN_2586; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2588 = 6'h13 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_19 : _GEN_2587; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2589 = 6'h14 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_20 : _GEN_2588; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2590 = 6'h15 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_21 : _GEN_2589; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2591 = 6'h16 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_22 : _GEN_2590; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2592 = 6'h17 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_23 : _GEN_2591; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2593 = 6'h18 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_24 : _GEN_2592; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2594 = 6'h19 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_25 : _GEN_2593; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2595 = 6'h1a == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_26 : _GEN_2594; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2596 = 6'h1b == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_27 : _GEN_2595; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2597 = 6'h1c == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_28 : _GEN_2596; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2598 = 6'h1d == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_29 : _GEN_2597; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2599 = 6'h1e == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_30 : _GEN_2598; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2600 = 6'h1f == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_31 : _GEN_2599; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2601 = 6'h20 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_32 : _GEN_2600; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2602 = 6'h21 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_33 : _GEN_2601; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2603 = 6'h22 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_34 : _GEN_2602; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2604 = 6'h23 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_35 : _GEN_2603; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2605 = 6'h24 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_36 : _GEN_2604; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2606 = 6'h25 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_37 : _GEN_2605; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2607 = 6'h26 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_38 : _GEN_2606; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2608 = 6'h27 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_39 : _GEN_2607; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2609 = 6'h28 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_40 : _GEN_2608; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2610 = 6'h29 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_41 : _GEN_2609; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2611 = 6'h2a == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_42 : _GEN_2610; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2612 = 6'h2b == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_43 : _GEN_2611; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2613 = 6'h2c == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_44 : _GEN_2612; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2614 = 6'h2d == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_45 : _GEN_2613; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2615 = 6'h2e == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_46 : _GEN_2614; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2616 = 6'h2f == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_47 : _GEN_2615; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2617 = 6'h30 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_48 : _GEN_2616; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2618 = 6'h31 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_49 : _GEN_2617; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2619 = 6'h32 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_50 : _GEN_2618; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2620 = 6'h33 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_51 : _GEN_2619; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2621 = 6'h34 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_52 : _GEN_2620; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2622 = 6'h35 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_53 : _GEN_2621; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2623 = 6'h36 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_54 : _GEN_2622; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2624 = 6'h37 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_55 : _GEN_2623; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2625 = 6'h38 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_56 : _GEN_2624; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2626 = 6'h39 == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_57 : _GEN_2625; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2627 = 6'h3a == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_58 : _GEN_2626; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2628 = 6'h3b == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_59 : _GEN_2627; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2629 = 6'h3c == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_60 : _GEN_2628; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2630 = 6'h3d == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_61 : _GEN_2629; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2631 = 6'h3e == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_62 : _GEN_2630; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_39 = 6'h3f == _myTriMemVec2_7_T_1[5:0] ? myHhdoutVec_63 : _GEN_2631; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2634 = 6'h1 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2635 = 6'h2 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_2 : _GEN_2634; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2636 = 6'h3 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_3 : _GEN_2635; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2637 = 6'h4 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_4 : _GEN_2636; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2638 = 6'h5 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_5 : _GEN_2637; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2639 = 6'h6 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_6 : _GEN_2638; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2640 = 6'h7 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_7 : _GEN_2639; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2641 = 6'h8 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_8 : _GEN_2640; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2642 = 6'h9 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_9 : _GEN_2641; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2643 = 6'ha == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_10 : _GEN_2642; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2644 = 6'hb == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_11 : _GEN_2643; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2645 = 6'hc == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_12 : _GEN_2644; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2646 = 6'hd == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_13 : _GEN_2645; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2647 = 6'he == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_14 : _GEN_2646; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2648 = 6'hf == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_15 : _GEN_2647; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2649 = 6'h10 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_16 : _GEN_2648; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2650 = 6'h11 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_17 : _GEN_2649; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2651 = 6'h12 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_18 : _GEN_2650; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2652 = 6'h13 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_19 : _GEN_2651; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2653 = 6'h14 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_20 : _GEN_2652; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2654 = 6'h15 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_21 : _GEN_2653; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2655 = 6'h16 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_22 : _GEN_2654; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2656 = 6'h17 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_23 : _GEN_2655; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2657 = 6'h18 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_24 : _GEN_2656; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2658 = 6'h19 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_25 : _GEN_2657; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2659 = 6'h1a == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_26 : _GEN_2658; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2660 = 6'h1b == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_27 : _GEN_2659; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2661 = 6'h1c == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_28 : _GEN_2660; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2662 = 6'h1d == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_29 : _GEN_2661; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2663 = 6'h1e == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_30 : _GEN_2662; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2664 = 6'h1f == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_31 : _GEN_2663; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2665 = 6'h20 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_32 : _GEN_2664; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2666 = 6'h21 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_33 : _GEN_2665; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2667 = 6'h22 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_34 : _GEN_2666; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2668 = 6'h23 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_35 : _GEN_2667; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2669 = 6'h24 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_36 : _GEN_2668; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2670 = 6'h25 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_37 : _GEN_2669; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2671 = 6'h26 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_38 : _GEN_2670; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2672 = 6'h27 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_39 : _GEN_2671; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2673 = 6'h28 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_40 : _GEN_2672; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2674 = 6'h29 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_41 : _GEN_2673; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2675 = 6'h2a == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_42 : _GEN_2674; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2676 = 6'h2b == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_43 : _GEN_2675; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2677 = 6'h2c == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_44 : _GEN_2676; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2678 = 6'h2d == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_45 : _GEN_2677; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2679 = 6'h2e == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_46 : _GEN_2678; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2680 = 6'h2f == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_47 : _GEN_2679; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2681 = 6'h30 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_48 : _GEN_2680; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2682 = 6'h31 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_49 : _GEN_2681; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2683 = 6'h32 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_50 : _GEN_2682; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2684 = 6'h33 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_51 : _GEN_2683; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2685 = 6'h34 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_52 : _GEN_2684; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2686 = 6'h35 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_53 : _GEN_2685; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2687 = 6'h36 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_54 : _GEN_2686; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2688 = 6'h37 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_55 : _GEN_2687; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2689 = 6'h38 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_56 : _GEN_2688; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2690 = 6'h39 == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_57 : _GEN_2689; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2691 = 6'h3a == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_58 : _GEN_2690; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2692 = 6'h3b == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_59 : _GEN_2691; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2693 = 6'h3c == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_60 : _GEN_2692; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2694 = 6'h3d == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_61 : _GEN_2693; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2695 = 6'h3e == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_62 : _GEN_2694; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_38 = 6'h3f == _myTriMemVec2_6_T_1[5:0] ? myHhdoutVec_63 : _GEN_2695; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2698 = 6'h1 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2699 = 6'h2 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_2 : _GEN_2698; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2700 = 6'h3 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_3 : _GEN_2699; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2701 = 6'h4 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_4 : _GEN_2700; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2702 = 6'h5 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_5 : _GEN_2701; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2703 = 6'h6 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_6 : _GEN_2702; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2704 = 6'h7 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_7 : _GEN_2703; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2705 = 6'h8 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_8 : _GEN_2704; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2706 = 6'h9 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_9 : _GEN_2705; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2707 = 6'ha == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_10 : _GEN_2706; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2708 = 6'hb == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_11 : _GEN_2707; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2709 = 6'hc == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_12 : _GEN_2708; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2710 = 6'hd == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_13 : _GEN_2709; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2711 = 6'he == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_14 : _GEN_2710; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2712 = 6'hf == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_15 : _GEN_2711; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2713 = 6'h10 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_16 : _GEN_2712; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2714 = 6'h11 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_17 : _GEN_2713; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2715 = 6'h12 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_18 : _GEN_2714; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2716 = 6'h13 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_19 : _GEN_2715; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2717 = 6'h14 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_20 : _GEN_2716; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2718 = 6'h15 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_21 : _GEN_2717; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2719 = 6'h16 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_22 : _GEN_2718; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2720 = 6'h17 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_23 : _GEN_2719; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2721 = 6'h18 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_24 : _GEN_2720; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2722 = 6'h19 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_25 : _GEN_2721; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2723 = 6'h1a == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_26 : _GEN_2722; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2724 = 6'h1b == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_27 : _GEN_2723; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2725 = 6'h1c == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_28 : _GEN_2724; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2726 = 6'h1d == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_29 : _GEN_2725; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2727 = 6'h1e == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_30 : _GEN_2726; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2728 = 6'h1f == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_31 : _GEN_2727; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2729 = 6'h20 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_32 : _GEN_2728; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2730 = 6'h21 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_33 : _GEN_2729; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2731 = 6'h22 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_34 : _GEN_2730; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2732 = 6'h23 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_35 : _GEN_2731; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2733 = 6'h24 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_36 : _GEN_2732; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2734 = 6'h25 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_37 : _GEN_2733; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2735 = 6'h26 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_38 : _GEN_2734; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2736 = 6'h27 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_39 : _GEN_2735; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2737 = 6'h28 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_40 : _GEN_2736; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2738 = 6'h29 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_41 : _GEN_2737; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2739 = 6'h2a == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_42 : _GEN_2738; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2740 = 6'h2b == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_43 : _GEN_2739; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2741 = 6'h2c == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_44 : _GEN_2740; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2742 = 6'h2d == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_45 : _GEN_2741; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2743 = 6'h2e == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_46 : _GEN_2742; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2744 = 6'h2f == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_47 : _GEN_2743; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2745 = 6'h30 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_48 : _GEN_2744; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2746 = 6'h31 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_49 : _GEN_2745; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2747 = 6'h32 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_50 : _GEN_2746; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2748 = 6'h33 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_51 : _GEN_2747; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2749 = 6'h34 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_52 : _GEN_2748; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2750 = 6'h35 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_53 : _GEN_2749; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2751 = 6'h36 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_54 : _GEN_2750; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2752 = 6'h37 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_55 : _GEN_2751; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2753 = 6'h38 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_56 : _GEN_2752; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2754 = 6'h39 == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_57 : _GEN_2753; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2755 = 6'h3a == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_58 : _GEN_2754; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2756 = 6'h3b == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_59 : _GEN_2755; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2757 = 6'h3c == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_60 : _GEN_2756; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2758 = 6'h3d == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_61 : _GEN_2757; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2759 = 6'h3e == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_62 : _GEN_2758; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_37 = 6'h3f == _myTriMemVec2_5_T_1[5:0] ? myHhdoutVec_63 : _GEN_2759; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2762 = 6'h1 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2763 = 6'h2 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_2 : _GEN_2762; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2764 = 6'h3 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_3 : _GEN_2763; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2765 = 6'h4 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_4 : _GEN_2764; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2766 = 6'h5 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_5 : _GEN_2765; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2767 = 6'h6 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_6 : _GEN_2766; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2768 = 6'h7 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_7 : _GEN_2767; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2769 = 6'h8 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_8 : _GEN_2768; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2770 = 6'h9 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_9 : _GEN_2769; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2771 = 6'ha == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_10 : _GEN_2770; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2772 = 6'hb == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_11 : _GEN_2771; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2773 = 6'hc == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_12 : _GEN_2772; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2774 = 6'hd == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_13 : _GEN_2773; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2775 = 6'he == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_14 : _GEN_2774; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2776 = 6'hf == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_15 : _GEN_2775; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2777 = 6'h10 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_16 : _GEN_2776; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2778 = 6'h11 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_17 : _GEN_2777; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2779 = 6'h12 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_18 : _GEN_2778; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2780 = 6'h13 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_19 : _GEN_2779; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2781 = 6'h14 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_20 : _GEN_2780; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2782 = 6'h15 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_21 : _GEN_2781; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2783 = 6'h16 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_22 : _GEN_2782; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2784 = 6'h17 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_23 : _GEN_2783; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2785 = 6'h18 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_24 : _GEN_2784; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2786 = 6'h19 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_25 : _GEN_2785; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2787 = 6'h1a == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_26 : _GEN_2786; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2788 = 6'h1b == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_27 : _GEN_2787; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2789 = 6'h1c == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_28 : _GEN_2788; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2790 = 6'h1d == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_29 : _GEN_2789; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2791 = 6'h1e == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_30 : _GEN_2790; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2792 = 6'h1f == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_31 : _GEN_2791; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2793 = 6'h20 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_32 : _GEN_2792; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2794 = 6'h21 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_33 : _GEN_2793; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2795 = 6'h22 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_34 : _GEN_2794; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2796 = 6'h23 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_35 : _GEN_2795; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2797 = 6'h24 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_36 : _GEN_2796; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2798 = 6'h25 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_37 : _GEN_2797; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2799 = 6'h26 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_38 : _GEN_2798; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2800 = 6'h27 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_39 : _GEN_2799; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2801 = 6'h28 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_40 : _GEN_2800; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2802 = 6'h29 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_41 : _GEN_2801; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2803 = 6'h2a == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_42 : _GEN_2802; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2804 = 6'h2b == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_43 : _GEN_2803; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2805 = 6'h2c == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_44 : _GEN_2804; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2806 = 6'h2d == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_45 : _GEN_2805; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2807 = 6'h2e == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_46 : _GEN_2806; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2808 = 6'h2f == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_47 : _GEN_2807; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2809 = 6'h30 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_48 : _GEN_2808; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2810 = 6'h31 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_49 : _GEN_2809; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2811 = 6'h32 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_50 : _GEN_2810; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2812 = 6'h33 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_51 : _GEN_2811; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2813 = 6'h34 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_52 : _GEN_2812; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2814 = 6'h35 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_53 : _GEN_2813; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2815 = 6'h36 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_54 : _GEN_2814; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2816 = 6'h37 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_55 : _GEN_2815; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2817 = 6'h38 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_56 : _GEN_2816; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2818 = 6'h39 == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_57 : _GEN_2817; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2819 = 6'h3a == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_58 : _GEN_2818; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2820 = 6'h3b == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_59 : _GEN_2819; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2821 = 6'h3c == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_60 : _GEN_2820; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2822 = 6'h3d == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_61 : _GEN_2821; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2823 = 6'h3e == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_62 : _GEN_2822; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_36 = 6'h3f == _myTriMemVec2_4_T_1[5:0] ? myHhdoutVec_63 : _GEN_2823; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2826 = 6'h1 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2827 = 6'h2 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_2 : _GEN_2826; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2828 = 6'h3 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_3 : _GEN_2827; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2829 = 6'h4 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_4 : _GEN_2828; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2830 = 6'h5 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_5 : _GEN_2829; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2831 = 6'h6 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_6 : _GEN_2830; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2832 = 6'h7 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_7 : _GEN_2831; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2833 = 6'h8 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_8 : _GEN_2832; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2834 = 6'h9 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_9 : _GEN_2833; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2835 = 6'ha == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_10 : _GEN_2834; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2836 = 6'hb == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_11 : _GEN_2835; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2837 = 6'hc == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_12 : _GEN_2836; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2838 = 6'hd == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_13 : _GEN_2837; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2839 = 6'he == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_14 : _GEN_2838; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2840 = 6'hf == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_15 : _GEN_2839; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2841 = 6'h10 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_16 : _GEN_2840; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2842 = 6'h11 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_17 : _GEN_2841; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2843 = 6'h12 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_18 : _GEN_2842; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2844 = 6'h13 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_19 : _GEN_2843; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2845 = 6'h14 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_20 : _GEN_2844; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2846 = 6'h15 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_21 : _GEN_2845; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2847 = 6'h16 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_22 : _GEN_2846; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2848 = 6'h17 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_23 : _GEN_2847; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2849 = 6'h18 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_24 : _GEN_2848; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2850 = 6'h19 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_25 : _GEN_2849; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2851 = 6'h1a == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_26 : _GEN_2850; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2852 = 6'h1b == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_27 : _GEN_2851; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2853 = 6'h1c == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_28 : _GEN_2852; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2854 = 6'h1d == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_29 : _GEN_2853; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2855 = 6'h1e == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_30 : _GEN_2854; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2856 = 6'h1f == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_31 : _GEN_2855; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2857 = 6'h20 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_32 : _GEN_2856; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2858 = 6'h21 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_33 : _GEN_2857; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2859 = 6'h22 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_34 : _GEN_2858; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2860 = 6'h23 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_35 : _GEN_2859; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2861 = 6'h24 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_36 : _GEN_2860; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2862 = 6'h25 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_37 : _GEN_2861; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2863 = 6'h26 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_38 : _GEN_2862; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2864 = 6'h27 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_39 : _GEN_2863; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2865 = 6'h28 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_40 : _GEN_2864; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2866 = 6'h29 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_41 : _GEN_2865; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2867 = 6'h2a == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_42 : _GEN_2866; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2868 = 6'h2b == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_43 : _GEN_2867; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2869 = 6'h2c == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_44 : _GEN_2868; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2870 = 6'h2d == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_45 : _GEN_2869; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2871 = 6'h2e == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_46 : _GEN_2870; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2872 = 6'h2f == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_47 : _GEN_2871; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2873 = 6'h30 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_48 : _GEN_2872; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2874 = 6'h31 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_49 : _GEN_2873; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2875 = 6'h32 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_50 : _GEN_2874; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2876 = 6'h33 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_51 : _GEN_2875; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2877 = 6'h34 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_52 : _GEN_2876; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2878 = 6'h35 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_53 : _GEN_2877; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2879 = 6'h36 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_54 : _GEN_2878; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2880 = 6'h37 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_55 : _GEN_2879; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2881 = 6'h38 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_56 : _GEN_2880; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2882 = 6'h39 == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_57 : _GEN_2881; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2883 = 6'h3a == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_58 : _GEN_2882; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2884 = 6'h3b == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_59 : _GEN_2883; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2885 = 6'h3c == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_60 : _GEN_2884; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2886 = 6'h3d == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_61 : _GEN_2885; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2887 = 6'h3e == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_62 : _GEN_2886; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_35 = 6'h3f == _myTriMemVec2_3_T_1[5:0] ? myHhdoutVec_63 : _GEN_2887; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2890 = 6'h1 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2891 = 6'h2 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_2 : _GEN_2890; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2892 = 6'h3 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_3 : _GEN_2891; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2893 = 6'h4 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_4 : _GEN_2892; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2894 = 6'h5 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_5 : _GEN_2893; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2895 = 6'h6 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_6 : _GEN_2894; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2896 = 6'h7 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_7 : _GEN_2895; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2897 = 6'h8 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_8 : _GEN_2896; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2898 = 6'h9 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_9 : _GEN_2897; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2899 = 6'ha == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_10 : _GEN_2898; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2900 = 6'hb == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_11 : _GEN_2899; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2901 = 6'hc == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_12 : _GEN_2900; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2902 = 6'hd == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_13 : _GEN_2901; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2903 = 6'he == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_14 : _GEN_2902; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2904 = 6'hf == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_15 : _GEN_2903; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2905 = 6'h10 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_16 : _GEN_2904; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2906 = 6'h11 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_17 : _GEN_2905; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2907 = 6'h12 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_18 : _GEN_2906; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2908 = 6'h13 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_19 : _GEN_2907; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2909 = 6'h14 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_20 : _GEN_2908; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2910 = 6'h15 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_21 : _GEN_2909; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2911 = 6'h16 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_22 : _GEN_2910; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2912 = 6'h17 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_23 : _GEN_2911; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2913 = 6'h18 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_24 : _GEN_2912; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2914 = 6'h19 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_25 : _GEN_2913; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2915 = 6'h1a == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_26 : _GEN_2914; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2916 = 6'h1b == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_27 : _GEN_2915; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2917 = 6'h1c == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_28 : _GEN_2916; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2918 = 6'h1d == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_29 : _GEN_2917; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2919 = 6'h1e == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_30 : _GEN_2918; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2920 = 6'h1f == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_31 : _GEN_2919; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2921 = 6'h20 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_32 : _GEN_2920; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2922 = 6'h21 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_33 : _GEN_2921; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2923 = 6'h22 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_34 : _GEN_2922; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2924 = 6'h23 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_35 : _GEN_2923; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2925 = 6'h24 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_36 : _GEN_2924; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2926 = 6'h25 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_37 : _GEN_2925; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2927 = 6'h26 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_38 : _GEN_2926; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2928 = 6'h27 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_39 : _GEN_2927; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2929 = 6'h28 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_40 : _GEN_2928; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2930 = 6'h29 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_41 : _GEN_2929; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2931 = 6'h2a == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_42 : _GEN_2930; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2932 = 6'h2b == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_43 : _GEN_2931; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2933 = 6'h2c == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_44 : _GEN_2932; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2934 = 6'h2d == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_45 : _GEN_2933; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2935 = 6'h2e == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_46 : _GEN_2934; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2936 = 6'h2f == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_47 : _GEN_2935; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2937 = 6'h30 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_48 : _GEN_2936; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2938 = 6'h31 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_49 : _GEN_2937; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2939 = 6'h32 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_50 : _GEN_2938; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2940 = 6'h33 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_51 : _GEN_2939; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2941 = 6'h34 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_52 : _GEN_2940; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2942 = 6'h35 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_53 : _GEN_2941; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2943 = 6'h36 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_54 : _GEN_2942; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2944 = 6'h37 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_55 : _GEN_2943; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2945 = 6'h38 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_56 : _GEN_2944; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2946 = 6'h39 == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_57 : _GEN_2945; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2947 = 6'h3a == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_58 : _GEN_2946; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2948 = 6'h3b == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_59 : _GEN_2947; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2949 = 6'h3c == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_60 : _GEN_2948; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2950 = 6'h3d == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_61 : _GEN_2949; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2951 = 6'h3e == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_62 : _GEN_2950; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_34 = 6'h3f == _myTriMemVec2_2_T_1[5:0] ? myHhdoutVec_63 : _GEN_2951; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2954 = 6'h1 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2955 = 6'h2 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_2 : _GEN_2954; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2956 = 6'h3 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_3 : _GEN_2955; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2957 = 6'h4 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_4 : _GEN_2956; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2958 = 6'h5 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_5 : _GEN_2957; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2959 = 6'h6 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_6 : _GEN_2958; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2960 = 6'h7 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_7 : _GEN_2959; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2961 = 6'h8 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_8 : _GEN_2960; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2962 = 6'h9 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_9 : _GEN_2961; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2963 = 6'ha == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_10 : _GEN_2962; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2964 = 6'hb == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_11 : _GEN_2963; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2965 = 6'hc == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_12 : _GEN_2964; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2966 = 6'hd == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_13 : _GEN_2965; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2967 = 6'he == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_14 : _GEN_2966; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2968 = 6'hf == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_15 : _GEN_2967; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2969 = 6'h10 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_16 : _GEN_2968; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2970 = 6'h11 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_17 : _GEN_2969; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2971 = 6'h12 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_18 : _GEN_2970; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2972 = 6'h13 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_19 : _GEN_2971; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2973 = 6'h14 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_20 : _GEN_2972; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2974 = 6'h15 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_21 : _GEN_2973; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2975 = 6'h16 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_22 : _GEN_2974; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2976 = 6'h17 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_23 : _GEN_2975; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2977 = 6'h18 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_24 : _GEN_2976; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2978 = 6'h19 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_25 : _GEN_2977; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2979 = 6'h1a == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_26 : _GEN_2978; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2980 = 6'h1b == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_27 : _GEN_2979; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2981 = 6'h1c == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_28 : _GEN_2980; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2982 = 6'h1d == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_29 : _GEN_2981; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2983 = 6'h1e == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_30 : _GEN_2982; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2984 = 6'h1f == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_31 : _GEN_2983; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2985 = 6'h20 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_32 : _GEN_2984; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2986 = 6'h21 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_33 : _GEN_2985; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2987 = 6'h22 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_34 : _GEN_2986; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2988 = 6'h23 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_35 : _GEN_2987; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2989 = 6'h24 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_36 : _GEN_2988; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2990 = 6'h25 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_37 : _GEN_2989; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2991 = 6'h26 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_38 : _GEN_2990; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2992 = 6'h27 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_39 : _GEN_2991; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2993 = 6'h28 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_40 : _GEN_2992; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2994 = 6'h29 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_41 : _GEN_2993; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2995 = 6'h2a == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_42 : _GEN_2994; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2996 = 6'h2b == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_43 : _GEN_2995; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2997 = 6'h2c == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_44 : _GEN_2996; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2998 = 6'h2d == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_45 : _GEN_2997; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_2999 = 6'h2e == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_46 : _GEN_2998; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3000 = 6'h2f == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_47 : _GEN_2999; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3001 = 6'h30 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_48 : _GEN_3000; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3002 = 6'h31 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_49 : _GEN_3001; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3003 = 6'h32 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_50 : _GEN_3002; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3004 = 6'h33 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_51 : _GEN_3003; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3005 = 6'h34 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_52 : _GEN_3004; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3006 = 6'h35 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_53 : _GEN_3005; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3007 = 6'h36 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_54 : _GEN_3006; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3008 = 6'h37 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_55 : _GEN_3007; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3009 = 6'h38 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_56 : _GEN_3008; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3010 = 6'h39 == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_57 : _GEN_3009; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3011 = 6'h3a == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_58 : _GEN_3010; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3012 = 6'h3b == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_59 : _GEN_3011; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3013 = 6'h3c == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_60 : _GEN_3012; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3014 = 6'h3d == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_61 : _GEN_3013; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3015 = 6'h3e == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_62 : _GEN_3014; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_33 = 6'h3f == _myTriMemVec2_1_T_1[5:0] ? myHhdoutVec_63 : _GEN_3015; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3018 = 6'h1 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3019 = 6'h2 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_2 : _GEN_3018; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3020 = 6'h3 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_3 : _GEN_3019; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3021 = 6'h4 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_4 : _GEN_3020; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3022 = 6'h5 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_5 : _GEN_3021; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3023 = 6'h6 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_6 : _GEN_3022; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3024 = 6'h7 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_7 : _GEN_3023; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3025 = 6'h8 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_8 : _GEN_3024; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3026 = 6'h9 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_9 : _GEN_3025; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3027 = 6'ha == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_10 : _GEN_3026; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3028 = 6'hb == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_11 : _GEN_3027; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3029 = 6'hc == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_12 : _GEN_3028; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3030 = 6'hd == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_13 : _GEN_3029; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3031 = 6'he == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_14 : _GEN_3030; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3032 = 6'hf == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_15 : _GEN_3031; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3033 = 6'h10 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_16 : _GEN_3032; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3034 = 6'h11 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_17 : _GEN_3033; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3035 = 6'h12 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_18 : _GEN_3034; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3036 = 6'h13 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_19 : _GEN_3035; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3037 = 6'h14 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_20 : _GEN_3036; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3038 = 6'h15 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_21 : _GEN_3037; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3039 = 6'h16 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_22 : _GEN_3038; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3040 = 6'h17 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_23 : _GEN_3039; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3041 = 6'h18 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_24 : _GEN_3040; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3042 = 6'h19 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_25 : _GEN_3041; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3043 = 6'h1a == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_26 : _GEN_3042; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3044 = 6'h1b == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_27 : _GEN_3043; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3045 = 6'h1c == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_28 : _GEN_3044; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3046 = 6'h1d == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_29 : _GEN_3045; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3047 = 6'h1e == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_30 : _GEN_3046; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3048 = 6'h1f == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_31 : _GEN_3047; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3049 = 6'h20 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_32 : _GEN_3048; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3050 = 6'h21 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_33 : _GEN_3049; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3051 = 6'h22 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_34 : _GEN_3050; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3052 = 6'h23 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_35 : _GEN_3051; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3053 = 6'h24 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_36 : _GEN_3052; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3054 = 6'h25 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_37 : _GEN_3053; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3055 = 6'h26 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_38 : _GEN_3054; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3056 = 6'h27 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_39 : _GEN_3055; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3057 = 6'h28 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_40 : _GEN_3056; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3058 = 6'h29 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_41 : _GEN_3057; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3059 = 6'h2a == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_42 : _GEN_3058; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3060 = 6'h2b == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_43 : _GEN_3059; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3061 = 6'h2c == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_44 : _GEN_3060; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3062 = 6'h2d == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_45 : _GEN_3061; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3063 = 6'h2e == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_46 : _GEN_3062; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3064 = 6'h2f == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_47 : _GEN_3063; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3065 = 6'h30 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_48 : _GEN_3064; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3066 = 6'h31 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_49 : _GEN_3065; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3067 = 6'h32 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_50 : _GEN_3066; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3068 = 6'h33 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_51 : _GEN_3067; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3069 = 6'h34 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_52 : _GEN_3068; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3070 = 6'h35 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_53 : _GEN_3069; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3071 = 6'h36 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_54 : _GEN_3070; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3072 = 6'h37 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_55 : _GEN_3071; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3073 = 6'h38 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_56 : _GEN_3072; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3074 = 6'h39 == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_57 : _GEN_3073; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3075 = 6'h3a == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_58 : _GEN_3074; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3076 = 6'h3b == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_59 : _GEN_3075; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3077 = 6'h3c == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_60 : _GEN_3076; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3078 = 6'h3d == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_61 : _GEN_3077; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3079 = 6'h3e == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_62 : _GEN_3078; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_32 = 6'h3f == _myTriMemVec2_0_T_1[5:0] ? myHhdoutVec_63 : _GEN_3079; // @[hh_core.scala 149:{52,52}]
  wire [255:0] myHhdoutWire_hi_lo_lo = {myHhdoutVec2_39,myHhdoutVec2_38,myHhdoutVec2_37,myHhdoutVec2_36,myHhdoutVec2_35,
    myHhdoutVec2_34,myHhdoutVec2_33,myHhdoutVec2_32}; // @[hh_core.scala 153:42]
  wire [511:0] myHhdoutWire_hi_lo = {myHhdoutVec2_47,myHhdoutVec2_46,myHhdoutVec2_45,myHhdoutVec2_44,myHhdoutVec2_43,
    myHhdoutVec2_42,myHhdoutVec2_41,myHhdoutVec2_40,myHhdoutWire_hi_lo_lo}; // @[hh_core.scala 153:42]
  wire [1023:0] myHhdoutWire_hi = {myHhdoutVec2_63,myHhdoutVec2_62,myHhdoutVec2_61,myHhdoutVec2_60,myHhdoutVec2_59,
    myHhdoutVec2_58,myHhdoutVec2_57,myHhdoutVec2_56,myHhdoutWire_hi_hi_lo,myHhdoutWire_hi_lo}; // @[hh_core.scala 153:42]
  wire [15:0] _myHhdoutVec2_31_T_1 = 16'h20 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3082 = 6'h1 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3083 = 6'h2 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_2 : _GEN_3082; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3084 = 6'h3 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_3 : _GEN_3083; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3085 = 6'h4 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_4 : _GEN_3084; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3086 = 6'h5 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_5 : _GEN_3085; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3087 = 6'h6 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_6 : _GEN_3086; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3088 = 6'h7 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_7 : _GEN_3087; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3089 = 6'h8 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_8 : _GEN_3088; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3090 = 6'h9 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_9 : _GEN_3089; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3091 = 6'ha == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_10 : _GEN_3090; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3092 = 6'hb == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_11 : _GEN_3091; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3093 = 6'hc == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_12 : _GEN_3092; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3094 = 6'hd == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_13 : _GEN_3093; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3095 = 6'he == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_14 : _GEN_3094; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3096 = 6'hf == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_15 : _GEN_3095; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3097 = 6'h10 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_16 : _GEN_3096; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3098 = 6'h11 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_17 : _GEN_3097; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3099 = 6'h12 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_18 : _GEN_3098; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3100 = 6'h13 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_19 : _GEN_3099; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3101 = 6'h14 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_20 : _GEN_3100; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3102 = 6'h15 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_21 : _GEN_3101; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3103 = 6'h16 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_22 : _GEN_3102; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3104 = 6'h17 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_23 : _GEN_3103; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3105 = 6'h18 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_24 : _GEN_3104; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3106 = 6'h19 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_25 : _GEN_3105; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3107 = 6'h1a == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_26 : _GEN_3106; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3108 = 6'h1b == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_27 : _GEN_3107; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3109 = 6'h1c == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_28 : _GEN_3108; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3110 = 6'h1d == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_29 : _GEN_3109; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3111 = 6'h1e == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_30 : _GEN_3110; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3112 = 6'h1f == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_31 : _GEN_3111; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3113 = 6'h20 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_32 : _GEN_3112; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3114 = 6'h21 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_33 : _GEN_3113; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3115 = 6'h22 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_34 : _GEN_3114; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3116 = 6'h23 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_35 : _GEN_3115; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3117 = 6'h24 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_36 : _GEN_3116; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3118 = 6'h25 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_37 : _GEN_3117; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3119 = 6'h26 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_38 : _GEN_3118; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3120 = 6'h27 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_39 : _GEN_3119; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3121 = 6'h28 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_40 : _GEN_3120; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3122 = 6'h29 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_41 : _GEN_3121; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3123 = 6'h2a == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_42 : _GEN_3122; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3124 = 6'h2b == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_43 : _GEN_3123; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3125 = 6'h2c == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_44 : _GEN_3124; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3126 = 6'h2d == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_45 : _GEN_3125; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3127 = 6'h2e == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_46 : _GEN_3126; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3128 = 6'h2f == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_47 : _GEN_3127; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3129 = 6'h30 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_48 : _GEN_3128; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3130 = 6'h31 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_49 : _GEN_3129; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3131 = 6'h32 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_50 : _GEN_3130; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3132 = 6'h33 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_51 : _GEN_3131; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3133 = 6'h34 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_52 : _GEN_3132; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3134 = 6'h35 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_53 : _GEN_3133; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3135 = 6'h36 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_54 : _GEN_3134; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3136 = 6'h37 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_55 : _GEN_3135; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3137 = 6'h38 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_56 : _GEN_3136; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3138 = 6'h39 == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_57 : _GEN_3137; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3139 = 6'h3a == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_58 : _GEN_3138; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3140 = 6'h3b == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_59 : _GEN_3139; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3141 = 6'h3c == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_60 : _GEN_3140; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3142 = 6'h3d == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_61 : _GEN_3141; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3143 = 6'h3e == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_62 : _GEN_3142; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_31 = 6'h3f == _myHhdoutVec2_31_T_1[5:0] ? myHhdoutVec_63 : _GEN_3143; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_30_T_1 = 16'h21 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3146 = 6'h1 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3147 = 6'h2 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_2 : _GEN_3146; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3148 = 6'h3 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_3 : _GEN_3147; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3149 = 6'h4 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_4 : _GEN_3148; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3150 = 6'h5 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_5 : _GEN_3149; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3151 = 6'h6 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_6 : _GEN_3150; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3152 = 6'h7 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_7 : _GEN_3151; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3153 = 6'h8 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_8 : _GEN_3152; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3154 = 6'h9 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_9 : _GEN_3153; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3155 = 6'ha == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_10 : _GEN_3154; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3156 = 6'hb == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_11 : _GEN_3155; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3157 = 6'hc == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_12 : _GEN_3156; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3158 = 6'hd == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_13 : _GEN_3157; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3159 = 6'he == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_14 : _GEN_3158; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3160 = 6'hf == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_15 : _GEN_3159; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3161 = 6'h10 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_16 : _GEN_3160; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3162 = 6'h11 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_17 : _GEN_3161; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3163 = 6'h12 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_18 : _GEN_3162; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3164 = 6'h13 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_19 : _GEN_3163; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3165 = 6'h14 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_20 : _GEN_3164; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3166 = 6'h15 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_21 : _GEN_3165; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3167 = 6'h16 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_22 : _GEN_3166; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3168 = 6'h17 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_23 : _GEN_3167; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3169 = 6'h18 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_24 : _GEN_3168; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3170 = 6'h19 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_25 : _GEN_3169; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3171 = 6'h1a == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_26 : _GEN_3170; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3172 = 6'h1b == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_27 : _GEN_3171; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3173 = 6'h1c == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_28 : _GEN_3172; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3174 = 6'h1d == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_29 : _GEN_3173; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3175 = 6'h1e == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_30 : _GEN_3174; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3176 = 6'h1f == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_31 : _GEN_3175; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3177 = 6'h20 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_32 : _GEN_3176; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3178 = 6'h21 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_33 : _GEN_3177; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3179 = 6'h22 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_34 : _GEN_3178; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3180 = 6'h23 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_35 : _GEN_3179; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3181 = 6'h24 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_36 : _GEN_3180; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3182 = 6'h25 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_37 : _GEN_3181; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3183 = 6'h26 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_38 : _GEN_3182; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3184 = 6'h27 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_39 : _GEN_3183; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3185 = 6'h28 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_40 : _GEN_3184; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3186 = 6'h29 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_41 : _GEN_3185; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3187 = 6'h2a == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_42 : _GEN_3186; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3188 = 6'h2b == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_43 : _GEN_3187; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3189 = 6'h2c == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_44 : _GEN_3188; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3190 = 6'h2d == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_45 : _GEN_3189; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3191 = 6'h2e == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_46 : _GEN_3190; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3192 = 6'h2f == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_47 : _GEN_3191; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3193 = 6'h30 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_48 : _GEN_3192; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3194 = 6'h31 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_49 : _GEN_3193; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3195 = 6'h32 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_50 : _GEN_3194; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3196 = 6'h33 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_51 : _GEN_3195; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3197 = 6'h34 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_52 : _GEN_3196; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3198 = 6'h35 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_53 : _GEN_3197; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3199 = 6'h36 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_54 : _GEN_3198; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3200 = 6'h37 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_55 : _GEN_3199; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3201 = 6'h38 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_56 : _GEN_3200; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3202 = 6'h39 == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_57 : _GEN_3201; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3203 = 6'h3a == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_58 : _GEN_3202; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3204 = 6'h3b == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_59 : _GEN_3203; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3205 = 6'h3c == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_60 : _GEN_3204; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3206 = 6'h3d == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_61 : _GEN_3205; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3207 = 6'h3e == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_62 : _GEN_3206; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_30 = 6'h3f == _myHhdoutVec2_30_T_1[5:0] ? myHhdoutVec_63 : _GEN_3207; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_29_T_1 = 16'h22 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3210 = 6'h1 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3211 = 6'h2 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_2 : _GEN_3210; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3212 = 6'h3 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_3 : _GEN_3211; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3213 = 6'h4 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_4 : _GEN_3212; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3214 = 6'h5 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_5 : _GEN_3213; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3215 = 6'h6 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_6 : _GEN_3214; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3216 = 6'h7 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_7 : _GEN_3215; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3217 = 6'h8 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_8 : _GEN_3216; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3218 = 6'h9 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_9 : _GEN_3217; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3219 = 6'ha == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_10 : _GEN_3218; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3220 = 6'hb == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_11 : _GEN_3219; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3221 = 6'hc == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_12 : _GEN_3220; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3222 = 6'hd == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_13 : _GEN_3221; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3223 = 6'he == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_14 : _GEN_3222; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3224 = 6'hf == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_15 : _GEN_3223; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3225 = 6'h10 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_16 : _GEN_3224; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3226 = 6'h11 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_17 : _GEN_3225; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3227 = 6'h12 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_18 : _GEN_3226; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3228 = 6'h13 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_19 : _GEN_3227; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3229 = 6'h14 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_20 : _GEN_3228; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3230 = 6'h15 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_21 : _GEN_3229; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3231 = 6'h16 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_22 : _GEN_3230; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3232 = 6'h17 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_23 : _GEN_3231; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3233 = 6'h18 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_24 : _GEN_3232; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3234 = 6'h19 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_25 : _GEN_3233; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3235 = 6'h1a == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_26 : _GEN_3234; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3236 = 6'h1b == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_27 : _GEN_3235; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3237 = 6'h1c == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_28 : _GEN_3236; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3238 = 6'h1d == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_29 : _GEN_3237; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3239 = 6'h1e == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_30 : _GEN_3238; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3240 = 6'h1f == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_31 : _GEN_3239; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3241 = 6'h20 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_32 : _GEN_3240; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3242 = 6'h21 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_33 : _GEN_3241; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3243 = 6'h22 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_34 : _GEN_3242; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3244 = 6'h23 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_35 : _GEN_3243; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3245 = 6'h24 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_36 : _GEN_3244; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3246 = 6'h25 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_37 : _GEN_3245; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3247 = 6'h26 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_38 : _GEN_3246; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3248 = 6'h27 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_39 : _GEN_3247; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3249 = 6'h28 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_40 : _GEN_3248; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3250 = 6'h29 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_41 : _GEN_3249; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3251 = 6'h2a == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_42 : _GEN_3250; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3252 = 6'h2b == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_43 : _GEN_3251; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3253 = 6'h2c == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_44 : _GEN_3252; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3254 = 6'h2d == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_45 : _GEN_3253; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3255 = 6'h2e == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_46 : _GEN_3254; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3256 = 6'h2f == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_47 : _GEN_3255; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3257 = 6'h30 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_48 : _GEN_3256; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3258 = 6'h31 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_49 : _GEN_3257; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3259 = 6'h32 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_50 : _GEN_3258; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3260 = 6'h33 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_51 : _GEN_3259; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3261 = 6'h34 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_52 : _GEN_3260; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3262 = 6'h35 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_53 : _GEN_3261; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3263 = 6'h36 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_54 : _GEN_3262; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3264 = 6'h37 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_55 : _GEN_3263; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3265 = 6'h38 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_56 : _GEN_3264; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3266 = 6'h39 == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_57 : _GEN_3265; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3267 = 6'h3a == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_58 : _GEN_3266; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3268 = 6'h3b == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_59 : _GEN_3267; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3269 = 6'h3c == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_60 : _GEN_3268; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3270 = 6'h3d == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_61 : _GEN_3269; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3271 = 6'h3e == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_62 : _GEN_3270; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_29 = 6'h3f == _myHhdoutVec2_29_T_1[5:0] ? myHhdoutVec_63 : _GEN_3271; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_28_T_1 = 16'h23 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3274 = 6'h1 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3275 = 6'h2 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_2 : _GEN_3274; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3276 = 6'h3 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_3 : _GEN_3275; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3277 = 6'h4 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_4 : _GEN_3276; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3278 = 6'h5 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_5 : _GEN_3277; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3279 = 6'h6 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_6 : _GEN_3278; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3280 = 6'h7 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_7 : _GEN_3279; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3281 = 6'h8 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_8 : _GEN_3280; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3282 = 6'h9 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_9 : _GEN_3281; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3283 = 6'ha == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_10 : _GEN_3282; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3284 = 6'hb == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_11 : _GEN_3283; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3285 = 6'hc == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_12 : _GEN_3284; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3286 = 6'hd == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_13 : _GEN_3285; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3287 = 6'he == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_14 : _GEN_3286; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3288 = 6'hf == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_15 : _GEN_3287; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3289 = 6'h10 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_16 : _GEN_3288; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3290 = 6'h11 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_17 : _GEN_3289; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3291 = 6'h12 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_18 : _GEN_3290; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3292 = 6'h13 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_19 : _GEN_3291; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3293 = 6'h14 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_20 : _GEN_3292; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3294 = 6'h15 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_21 : _GEN_3293; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3295 = 6'h16 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_22 : _GEN_3294; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3296 = 6'h17 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_23 : _GEN_3295; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3297 = 6'h18 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_24 : _GEN_3296; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3298 = 6'h19 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_25 : _GEN_3297; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3299 = 6'h1a == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_26 : _GEN_3298; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3300 = 6'h1b == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_27 : _GEN_3299; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3301 = 6'h1c == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_28 : _GEN_3300; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3302 = 6'h1d == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_29 : _GEN_3301; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3303 = 6'h1e == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_30 : _GEN_3302; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3304 = 6'h1f == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_31 : _GEN_3303; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3305 = 6'h20 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_32 : _GEN_3304; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3306 = 6'h21 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_33 : _GEN_3305; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3307 = 6'h22 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_34 : _GEN_3306; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3308 = 6'h23 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_35 : _GEN_3307; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3309 = 6'h24 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_36 : _GEN_3308; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3310 = 6'h25 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_37 : _GEN_3309; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3311 = 6'h26 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_38 : _GEN_3310; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3312 = 6'h27 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_39 : _GEN_3311; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3313 = 6'h28 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_40 : _GEN_3312; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3314 = 6'h29 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_41 : _GEN_3313; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3315 = 6'h2a == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_42 : _GEN_3314; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3316 = 6'h2b == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_43 : _GEN_3315; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3317 = 6'h2c == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_44 : _GEN_3316; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3318 = 6'h2d == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_45 : _GEN_3317; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3319 = 6'h2e == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_46 : _GEN_3318; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3320 = 6'h2f == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_47 : _GEN_3319; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3321 = 6'h30 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_48 : _GEN_3320; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3322 = 6'h31 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_49 : _GEN_3321; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3323 = 6'h32 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_50 : _GEN_3322; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3324 = 6'h33 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_51 : _GEN_3323; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3325 = 6'h34 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_52 : _GEN_3324; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3326 = 6'h35 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_53 : _GEN_3325; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3327 = 6'h36 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_54 : _GEN_3326; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3328 = 6'h37 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_55 : _GEN_3327; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3329 = 6'h38 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_56 : _GEN_3328; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3330 = 6'h39 == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_57 : _GEN_3329; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3331 = 6'h3a == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_58 : _GEN_3330; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3332 = 6'h3b == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_59 : _GEN_3331; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3333 = 6'h3c == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_60 : _GEN_3332; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3334 = 6'h3d == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_61 : _GEN_3333; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3335 = 6'h3e == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_62 : _GEN_3334; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_28 = 6'h3f == _myHhdoutVec2_28_T_1[5:0] ? myHhdoutVec_63 : _GEN_3335; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_27_T_1 = 16'h24 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3338 = 6'h1 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3339 = 6'h2 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_2 : _GEN_3338; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3340 = 6'h3 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_3 : _GEN_3339; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3341 = 6'h4 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_4 : _GEN_3340; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3342 = 6'h5 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_5 : _GEN_3341; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3343 = 6'h6 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_6 : _GEN_3342; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3344 = 6'h7 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_7 : _GEN_3343; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3345 = 6'h8 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_8 : _GEN_3344; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3346 = 6'h9 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_9 : _GEN_3345; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3347 = 6'ha == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_10 : _GEN_3346; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3348 = 6'hb == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_11 : _GEN_3347; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3349 = 6'hc == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_12 : _GEN_3348; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3350 = 6'hd == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_13 : _GEN_3349; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3351 = 6'he == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_14 : _GEN_3350; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3352 = 6'hf == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_15 : _GEN_3351; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3353 = 6'h10 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_16 : _GEN_3352; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3354 = 6'h11 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_17 : _GEN_3353; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3355 = 6'h12 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_18 : _GEN_3354; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3356 = 6'h13 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_19 : _GEN_3355; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3357 = 6'h14 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_20 : _GEN_3356; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3358 = 6'h15 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_21 : _GEN_3357; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3359 = 6'h16 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_22 : _GEN_3358; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3360 = 6'h17 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_23 : _GEN_3359; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3361 = 6'h18 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_24 : _GEN_3360; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3362 = 6'h19 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_25 : _GEN_3361; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3363 = 6'h1a == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_26 : _GEN_3362; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3364 = 6'h1b == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_27 : _GEN_3363; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3365 = 6'h1c == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_28 : _GEN_3364; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3366 = 6'h1d == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_29 : _GEN_3365; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3367 = 6'h1e == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_30 : _GEN_3366; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3368 = 6'h1f == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_31 : _GEN_3367; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3369 = 6'h20 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_32 : _GEN_3368; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3370 = 6'h21 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_33 : _GEN_3369; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3371 = 6'h22 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_34 : _GEN_3370; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3372 = 6'h23 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_35 : _GEN_3371; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3373 = 6'h24 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_36 : _GEN_3372; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3374 = 6'h25 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_37 : _GEN_3373; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3375 = 6'h26 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_38 : _GEN_3374; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3376 = 6'h27 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_39 : _GEN_3375; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3377 = 6'h28 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_40 : _GEN_3376; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3378 = 6'h29 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_41 : _GEN_3377; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3379 = 6'h2a == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_42 : _GEN_3378; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3380 = 6'h2b == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_43 : _GEN_3379; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3381 = 6'h2c == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_44 : _GEN_3380; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3382 = 6'h2d == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_45 : _GEN_3381; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3383 = 6'h2e == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_46 : _GEN_3382; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3384 = 6'h2f == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_47 : _GEN_3383; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3385 = 6'h30 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_48 : _GEN_3384; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3386 = 6'h31 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_49 : _GEN_3385; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3387 = 6'h32 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_50 : _GEN_3386; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3388 = 6'h33 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_51 : _GEN_3387; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3389 = 6'h34 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_52 : _GEN_3388; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3390 = 6'h35 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_53 : _GEN_3389; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3391 = 6'h36 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_54 : _GEN_3390; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3392 = 6'h37 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_55 : _GEN_3391; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3393 = 6'h38 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_56 : _GEN_3392; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3394 = 6'h39 == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_57 : _GEN_3393; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3395 = 6'h3a == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_58 : _GEN_3394; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3396 = 6'h3b == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_59 : _GEN_3395; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3397 = 6'h3c == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_60 : _GEN_3396; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3398 = 6'h3d == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_61 : _GEN_3397; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3399 = 6'h3e == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_62 : _GEN_3398; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_27 = 6'h3f == _myHhdoutVec2_27_T_1[5:0] ? myHhdoutVec_63 : _GEN_3399; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_26_T_1 = 16'h25 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3402 = 6'h1 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3403 = 6'h2 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_2 : _GEN_3402; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3404 = 6'h3 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_3 : _GEN_3403; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3405 = 6'h4 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_4 : _GEN_3404; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3406 = 6'h5 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_5 : _GEN_3405; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3407 = 6'h6 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_6 : _GEN_3406; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3408 = 6'h7 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_7 : _GEN_3407; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3409 = 6'h8 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_8 : _GEN_3408; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3410 = 6'h9 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_9 : _GEN_3409; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3411 = 6'ha == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_10 : _GEN_3410; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3412 = 6'hb == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_11 : _GEN_3411; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3413 = 6'hc == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_12 : _GEN_3412; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3414 = 6'hd == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_13 : _GEN_3413; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3415 = 6'he == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_14 : _GEN_3414; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3416 = 6'hf == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_15 : _GEN_3415; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3417 = 6'h10 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_16 : _GEN_3416; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3418 = 6'h11 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_17 : _GEN_3417; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3419 = 6'h12 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_18 : _GEN_3418; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3420 = 6'h13 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_19 : _GEN_3419; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3421 = 6'h14 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_20 : _GEN_3420; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3422 = 6'h15 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_21 : _GEN_3421; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3423 = 6'h16 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_22 : _GEN_3422; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3424 = 6'h17 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_23 : _GEN_3423; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3425 = 6'h18 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_24 : _GEN_3424; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3426 = 6'h19 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_25 : _GEN_3425; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3427 = 6'h1a == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_26 : _GEN_3426; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3428 = 6'h1b == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_27 : _GEN_3427; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3429 = 6'h1c == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_28 : _GEN_3428; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3430 = 6'h1d == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_29 : _GEN_3429; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3431 = 6'h1e == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_30 : _GEN_3430; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3432 = 6'h1f == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_31 : _GEN_3431; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3433 = 6'h20 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_32 : _GEN_3432; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3434 = 6'h21 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_33 : _GEN_3433; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3435 = 6'h22 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_34 : _GEN_3434; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3436 = 6'h23 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_35 : _GEN_3435; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3437 = 6'h24 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_36 : _GEN_3436; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3438 = 6'h25 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_37 : _GEN_3437; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3439 = 6'h26 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_38 : _GEN_3438; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3440 = 6'h27 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_39 : _GEN_3439; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3441 = 6'h28 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_40 : _GEN_3440; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3442 = 6'h29 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_41 : _GEN_3441; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3443 = 6'h2a == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_42 : _GEN_3442; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3444 = 6'h2b == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_43 : _GEN_3443; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3445 = 6'h2c == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_44 : _GEN_3444; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3446 = 6'h2d == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_45 : _GEN_3445; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3447 = 6'h2e == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_46 : _GEN_3446; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3448 = 6'h2f == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_47 : _GEN_3447; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3449 = 6'h30 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_48 : _GEN_3448; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3450 = 6'h31 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_49 : _GEN_3449; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3451 = 6'h32 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_50 : _GEN_3450; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3452 = 6'h33 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_51 : _GEN_3451; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3453 = 6'h34 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_52 : _GEN_3452; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3454 = 6'h35 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_53 : _GEN_3453; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3455 = 6'h36 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_54 : _GEN_3454; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3456 = 6'h37 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_55 : _GEN_3455; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3457 = 6'h38 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_56 : _GEN_3456; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3458 = 6'h39 == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_57 : _GEN_3457; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3459 = 6'h3a == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_58 : _GEN_3458; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3460 = 6'h3b == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_59 : _GEN_3459; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3461 = 6'h3c == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_60 : _GEN_3460; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3462 = 6'h3d == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_61 : _GEN_3461; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3463 = 6'h3e == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_62 : _GEN_3462; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_26 = 6'h3f == _myHhdoutVec2_26_T_1[5:0] ? myHhdoutVec_63 : _GEN_3463; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_25_T_1 = 16'h26 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3466 = 6'h1 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3467 = 6'h2 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_2 : _GEN_3466; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3468 = 6'h3 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_3 : _GEN_3467; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3469 = 6'h4 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_4 : _GEN_3468; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3470 = 6'h5 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_5 : _GEN_3469; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3471 = 6'h6 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_6 : _GEN_3470; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3472 = 6'h7 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_7 : _GEN_3471; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3473 = 6'h8 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_8 : _GEN_3472; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3474 = 6'h9 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_9 : _GEN_3473; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3475 = 6'ha == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_10 : _GEN_3474; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3476 = 6'hb == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_11 : _GEN_3475; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3477 = 6'hc == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_12 : _GEN_3476; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3478 = 6'hd == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_13 : _GEN_3477; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3479 = 6'he == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_14 : _GEN_3478; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3480 = 6'hf == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_15 : _GEN_3479; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3481 = 6'h10 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_16 : _GEN_3480; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3482 = 6'h11 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_17 : _GEN_3481; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3483 = 6'h12 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_18 : _GEN_3482; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3484 = 6'h13 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_19 : _GEN_3483; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3485 = 6'h14 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_20 : _GEN_3484; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3486 = 6'h15 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_21 : _GEN_3485; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3487 = 6'h16 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_22 : _GEN_3486; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3488 = 6'h17 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_23 : _GEN_3487; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3489 = 6'h18 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_24 : _GEN_3488; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3490 = 6'h19 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_25 : _GEN_3489; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3491 = 6'h1a == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_26 : _GEN_3490; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3492 = 6'h1b == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_27 : _GEN_3491; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3493 = 6'h1c == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_28 : _GEN_3492; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3494 = 6'h1d == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_29 : _GEN_3493; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3495 = 6'h1e == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_30 : _GEN_3494; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3496 = 6'h1f == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_31 : _GEN_3495; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3497 = 6'h20 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_32 : _GEN_3496; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3498 = 6'h21 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_33 : _GEN_3497; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3499 = 6'h22 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_34 : _GEN_3498; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3500 = 6'h23 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_35 : _GEN_3499; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3501 = 6'h24 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_36 : _GEN_3500; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3502 = 6'h25 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_37 : _GEN_3501; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3503 = 6'h26 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_38 : _GEN_3502; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3504 = 6'h27 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_39 : _GEN_3503; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3505 = 6'h28 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_40 : _GEN_3504; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3506 = 6'h29 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_41 : _GEN_3505; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3507 = 6'h2a == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_42 : _GEN_3506; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3508 = 6'h2b == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_43 : _GEN_3507; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3509 = 6'h2c == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_44 : _GEN_3508; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3510 = 6'h2d == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_45 : _GEN_3509; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3511 = 6'h2e == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_46 : _GEN_3510; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3512 = 6'h2f == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_47 : _GEN_3511; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3513 = 6'h30 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_48 : _GEN_3512; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3514 = 6'h31 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_49 : _GEN_3513; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3515 = 6'h32 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_50 : _GEN_3514; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3516 = 6'h33 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_51 : _GEN_3515; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3517 = 6'h34 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_52 : _GEN_3516; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3518 = 6'h35 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_53 : _GEN_3517; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3519 = 6'h36 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_54 : _GEN_3518; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3520 = 6'h37 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_55 : _GEN_3519; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3521 = 6'h38 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_56 : _GEN_3520; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3522 = 6'h39 == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_57 : _GEN_3521; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3523 = 6'h3a == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_58 : _GEN_3522; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3524 = 6'h3b == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_59 : _GEN_3523; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3525 = 6'h3c == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_60 : _GEN_3524; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3526 = 6'h3d == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_61 : _GEN_3525; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3527 = 6'h3e == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_62 : _GEN_3526; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_25 = 6'h3f == _myHhdoutVec2_25_T_1[5:0] ? myHhdoutVec_63 : _GEN_3527; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_24_T_1 = 16'h27 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3530 = 6'h1 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3531 = 6'h2 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_2 : _GEN_3530; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3532 = 6'h3 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_3 : _GEN_3531; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3533 = 6'h4 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_4 : _GEN_3532; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3534 = 6'h5 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_5 : _GEN_3533; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3535 = 6'h6 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_6 : _GEN_3534; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3536 = 6'h7 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_7 : _GEN_3535; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3537 = 6'h8 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_8 : _GEN_3536; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3538 = 6'h9 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_9 : _GEN_3537; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3539 = 6'ha == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_10 : _GEN_3538; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3540 = 6'hb == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_11 : _GEN_3539; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3541 = 6'hc == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_12 : _GEN_3540; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3542 = 6'hd == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_13 : _GEN_3541; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3543 = 6'he == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_14 : _GEN_3542; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3544 = 6'hf == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_15 : _GEN_3543; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3545 = 6'h10 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_16 : _GEN_3544; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3546 = 6'h11 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_17 : _GEN_3545; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3547 = 6'h12 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_18 : _GEN_3546; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3548 = 6'h13 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_19 : _GEN_3547; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3549 = 6'h14 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_20 : _GEN_3548; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3550 = 6'h15 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_21 : _GEN_3549; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3551 = 6'h16 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_22 : _GEN_3550; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3552 = 6'h17 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_23 : _GEN_3551; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3553 = 6'h18 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_24 : _GEN_3552; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3554 = 6'h19 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_25 : _GEN_3553; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3555 = 6'h1a == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_26 : _GEN_3554; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3556 = 6'h1b == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_27 : _GEN_3555; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3557 = 6'h1c == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_28 : _GEN_3556; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3558 = 6'h1d == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_29 : _GEN_3557; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3559 = 6'h1e == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_30 : _GEN_3558; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3560 = 6'h1f == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_31 : _GEN_3559; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3561 = 6'h20 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_32 : _GEN_3560; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3562 = 6'h21 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_33 : _GEN_3561; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3563 = 6'h22 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_34 : _GEN_3562; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3564 = 6'h23 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_35 : _GEN_3563; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3565 = 6'h24 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_36 : _GEN_3564; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3566 = 6'h25 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_37 : _GEN_3565; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3567 = 6'h26 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_38 : _GEN_3566; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3568 = 6'h27 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_39 : _GEN_3567; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3569 = 6'h28 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_40 : _GEN_3568; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3570 = 6'h29 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_41 : _GEN_3569; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3571 = 6'h2a == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_42 : _GEN_3570; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3572 = 6'h2b == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_43 : _GEN_3571; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3573 = 6'h2c == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_44 : _GEN_3572; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3574 = 6'h2d == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_45 : _GEN_3573; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3575 = 6'h2e == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_46 : _GEN_3574; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3576 = 6'h2f == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_47 : _GEN_3575; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3577 = 6'h30 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_48 : _GEN_3576; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3578 = 6'h31 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_49 : _GEN_3577; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3579 = 6'h32 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_50 : _GEN_3578; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3580 = 6'h33 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_51 : _GEN_3579; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3581 = 6'h34 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_52 : _GEN_3580; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3582 = 6'h35 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_53 : _GEN_3581; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3583 = 6'h36 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_54 : _GEN_3582; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3584 = 6'h37 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_55 : _GEN_3583; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3585 = 6'h38 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_56 : _GEN_3584; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3586 = 6'h39 == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_57 : _GEN_3585; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3587 = 6'h3a == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_58 : _GEN_3586; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3588 = 6'h3b == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_59 : _GEN_3587; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3589 = 6'h3c == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_60 : _GEN_3588; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3590 = 6'h3d == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_61 : _GEN_3589; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3591 = 6'h3e == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_62 : _GEN_3590; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_24 = 6'h3f == _myHhdoutVec2_24_T_1[5:0] ? myHhdoutVec_63 : _GEN_3591; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_23_T_1 = 16'h28 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3594 = 6'h1 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3595 = 6'h2 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_2 : _GEN_3594; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3596 = 6'h3 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_3 : _GEN_3595; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3597 = 6'h4 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_4 : _GEN_3596; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3598 = 6'h5 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_5 : _GEN_3597; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3599 = 6'h6 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_6 : _GEN_3598; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3600 = 6'h7 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_7 : _GEN_3599; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3601 = 6'h8 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_8 : _GEN_3600; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3602 = 6'h9 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_9 : _GEN_3601; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3603 = 6'ha == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_10 : _GEN_3602; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3604 = 6'hb == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_11 : _GEN_3603; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3605 = 6'hc == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_12 : _GEN_3604; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3606 = 6'hd == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_13 : _GEN_3605; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3607 = 6'he == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_14 : _GEN_3606; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3608 = 6'hf == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_15 : _GEN_3607; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3609 = 6'h10 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_16 : _GEN_3608; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3610 = 6'h11 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_17 : _GEN_3609; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3611 = 6'h12 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_18 : _GEN_3610; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3612 = 6'h13 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_19 : _GEN_3611; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3613 = 6'h14 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_20 : _GEN_3612; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3614 = 6'h15 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_21 : _GEN_3613; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3615 = 6'h16 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_22 : _GEN_3614; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3616 = 6'h17 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_23 : _GEN_3615; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3617 = 6'h18 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_24 : _GEN_3616; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3618 = 6'h19 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_25 : _GEN_3617; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3619 = 6'h1a == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_26 : _GEN_3618; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3620 = 6'h1b == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_27 : _GEN_3619; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3621 = 6'h1c == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_28 : _GEN_3620; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3622 = 6'h1d == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_29 : _GEN_3621; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3623 = 6'h1e == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_30 : _GEN_3622; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3624 = 6'h1f == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_31 : _GEN_3623; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3625 = 6'h20 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_32 : _GEN_3624; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3626 = 6'h21 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_33 : _GEN_3625; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3627 = 6'h22 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_34 : _GEN_3626; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3628 = 6'h23 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_35 : _GEN_3627; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3629 = 6'h24 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_36 : _GEN_3628; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3630 = 6'h25 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_37 : _GEN_3629; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3631 = 6'h26 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_38 : _GEN_3630; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3632 = 6'h27 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_39 : _GEN_3631; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3633 = 6'h28 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_40 : _GEN_3632; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3634 = 6'h29 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_41 : _GEN_3633; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3635 = 6'h2a == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_42 : _GEN_3634; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3636 = 6'h2b == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_43 : _GEN_3635; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3637 = 6'h2c == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_44 : _GEN_3636; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3638 = 6'h2d == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_45 : _GEN_3637; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3639 = 6'h2e == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_46 : _GEN_3638; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3640 = 6'h2f == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_47 : _GEN_3639; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3641 = 6'h30 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_48 : _GEN_3640; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3642 = 6'h31 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_49 : _GEN_3641; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3643 = 6'h32 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_50 : _GEN_3642; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3644 = 6'h33 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_51 : _GEN_3643; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3645 = 6'h34 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_52 : _GEN_3644; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3646 = 6'h35 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_53 : _GEN_3645; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3647 = 6'h36 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_54 : _GEN_3646; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3648 = 6'h37 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_55 : _GEN_3647; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3649 = 6'h38 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_56 : _GEN_3648; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3650 = 6'h39 == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_57 : _GEN_3649; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3651 = 6'h3a == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_58 : _GEN_3650; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3652 = 6'h3b == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_59 : _GEN_3651; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3653 = 6'h3c == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_60 : _GEN_3652; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3654 = 6'h3d == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_61 : _GEN_3653; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3655 = 6'h3e == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_62 : _GEN_3654; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_23 = 6'h3f == _myHhdoutVec2_23_T_1[5:0] ? myHhdoutVec_63 : _GEN_3655; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_22_T_1 = 16'h29 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3658 = 6'h1 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3659 = 6'h2 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_2 : _GEN_3658; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3660 = 6'h3 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_3 : _GEN_3659; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3661 = 6'h4 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_4 : _GEN_3660; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3662 = 6'h5 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_5 : _GEN_3661; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3663 = 6'h6 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_6 : _GEN_3662; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3664 = 6'h7 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_7 : _GEN_3663; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3665 = 6'h8 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_8 : _GEN_3664; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3666 = 6'h9 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_9 : _GEN_3665; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3667 = 6'ha == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_10 : _GEN_3666; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3668 = 6'hb == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_11 : _GEN_3667; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3669 = 6'hc == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_12 : _GEN_3668; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3670 = 6'hd == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_13 : _GEN_3669; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3671 = 6'he == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_14 : _GEN_3670; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3672 = 6'hf == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_15 : _GEN_3671; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3673 = 6'h10 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_16 : _GEN_3672; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3674 = 6'h11 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_17 : _GEN_3673; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3675 = 6'h12 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_18 : _GEN_3674; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3676 = 6'h13 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_19 : _GEN_3675; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3677 = 6'h14 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_20 : _GEN_3676; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3678 = 6'h15 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_21 : _GEN_3677; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3679 = 6'h16 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_22 : _GEN_3678; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3680 = 6'h17 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_23 : _GEN_3679; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3681 = 6'h18 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_24 : _GEN_3680; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3682 = 6'h19 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_25 : _GEN_3681; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3683 = 6'h1a == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_26 : _GEN_3682; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3684 = 6'h1b == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_27 : _GEN_3683; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3685 = 6'h1c == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_28 : _GEN_3684; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3686 = 6'h1d == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_29 : _GEN_3685; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3687 = 6'h1e == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_30 : _GEN_3686; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3688 = 6'h1f == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_31 : _GEN_3687; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3689 = 6'h20 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_32 : _GEN_3688; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3690 = 6'h21 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_33 : _GEN_3689; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3691 = 6'h22 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_34 : _GEN_3690; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3692 = 6'h23 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_35 : _GEN_3691; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3693 = 6'h24 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_36 : _GEN_3692; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3694 = 6'h25 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_37 : _GEN_3693; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3695 = 6'h26 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_38 : _GEN_3694; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3696 = 6'h27 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_39 : _GEN_3695; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3697 = 6'h28 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_40 : _GEN_3696; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3698 = 6'h29 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_41 : _GEN_3697; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3699 = 6'h2a == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_42 : _GEN_3698; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3700 = 6'h2b == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_43 : _GEN_3699; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3701 = 6'h2c == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_44 : _GEN_3700; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3702 = 6'h2d == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_45 : _GEN_3701; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3703 = 6'h2e == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_46 : _GEN_3702; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3704 = 6'h2f == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_47 : _GEN_3703; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3705 = 6'h30 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_48 : _GEN_3704; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3706 = 6'h31 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_49 : _GEN_3705; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3707 = 6'h32 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_50 : _GEN_3706; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3708 = 6'h33 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_51 : _GEN_3707; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3709 = 6'h34 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_52 : _GEN_3708; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3710 = 6'h35 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_53 : _GEN_3709; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3711 = 6'h36 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_54 : _GEN_3710; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3712 = 6'h37 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_55 : _GEN_3711; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3713 = 6'h38 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_56 : _GEN_3712; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3714 = 6'h39 == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_57 : _GEN_3713; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3715 = 6'h3a == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_58 : _GEN_3714; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3716 = 6'h3b == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_59 : _GEN_3715; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3717 = 6'h3c == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_60 : _GEN_3716; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3718 = 6'h3d == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_61 : _GEN_3717; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3719 = 6'h3e == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_62 : _GEN_3718; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_22 = 6'h3f == _myHhdoutVec2_22_T_1[5:0] ? myHhdoutVec_63 : _GEN_3719; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_21_T_1 = 16'h2a + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3722 = 6'h1 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3723 = 6'h2 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_2 : _GEN_3722; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3724 = 6'h3 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_3 : _GEN_3723; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3725 = 6'h4 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_4 : _GEN_3724; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3726 = 6'h5 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_5 : _GEN_3725; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3727 = 6'h6 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_6 : _GEN_3726; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3728 = 6'h7 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_7 : _GEN_3727; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3729 = 6'h8 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_8 : _GEN_3728; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3730 = 6'h9 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_9 : _GEN_3729; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3731 = 6'ha == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_10 : _GEN_3730; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3732 = 6'hb == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_11 : _GEN_3731; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3733 = 6'hc == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_12 : _GEN_3732; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3734 = 6'hd == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_13 : _GEN_3733; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3735 = 6'he == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_14 : _GEN_3734; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3736 = 6'hf == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_15 : _GEN_3735; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3737 = 6'h10 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_16 : _GEN_3736; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3738 = 6'h11 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_17 : _GEN_3737; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3739 = 6'h12 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_18 : _GEN_3738; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3740 = 6'h13 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_19 : _GEN_3739; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3741 = 6'h14 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_20 : _GEN_3740; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3742 = 6'h15 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_21 : _GEN_3741; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3743 = 6'h16 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_22 : _GEN_3742; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3744 = 6'h17 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_23 : _GEN_3743; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3745 = 6'h18 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_24 : _GEN_3744; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3746 = 6'h19 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_25 : _GEN_3745; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3747 = 6'h1a == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_26 : _GEN_3746; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3748 = 6'h1b == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_27 : _GEN_3747; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3749 = 6'h1c == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_28 : _GEN_3748; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3750 = 6'h1d == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_29 : _GEN_3749; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3751 = 6'h1e == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_30 : _GEN_3750; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3752 = 6'h1f == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_31 : _GEN_3751; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3753 = 6'h20 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_32 : _GEN_3752; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3754 = 6'h21 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_33 : _GEN_3753; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3755 = 6'h22 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_34 : _GEN_3754; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3756 = 6'h23 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_35 : _GEN_3755; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3757 = 6'h24 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_36 : _GEN_3756; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3758 = 6'h25 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_37 : _GEN_3757; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3759 = 6'h26 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_38 : _GEN_3758; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3760 = 6'h27 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_39 : _GEN_3759; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3761 = 6'h28 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_40 : _GEN_3760; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3762 = 6'h29 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_41 : _GEN_3761; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3763 = 6'h2a == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_42 : _GEN_3762; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3764 = 6'h2b == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_43 : _GEN_3763; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3765 = 6'h2c == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_44 : _GEN_3764; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3766 = 6'h2d == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_45 : _GEN_3765; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3767 = 6'h2e == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_46 : _GEN_3766; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3768 = 6'h2f == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_47 : _GEN_3767; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3769 = 6'h30 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_48 : _GEN_3768; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3770 = 6'h31 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_49 : _GEN_3769; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3771 = 6'h32 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_50 : _GEN_3770; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3772 = 6'h33 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_51 : _GEN_3771; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3773 = 6'h34 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_52 : _GEN_3772; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3774 = 6'h35 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_53 : _GEN_3773; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3775 = 6'h36 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_54 : _GEN_3774; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3776 = 6'h37 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_55 : _GEN_3775; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3777 = 6'h38 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_56 : _GEN_3776; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3778 = 6'h39 == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_57 : _GEN_3777; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3779 = 6'h3a == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_58 : _GEN_3778; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3780 = 6'h3b == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_59 : _GEN_3779; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3781 = 6'h3c == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_60 : _GEN_3780; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3782 = 6'h3d == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_61 : _GEN_3781; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3783 = 6'h3e == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_62 : _GEN_3782; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_21 = 6'h3f == _myHhdoutVec2_21_T_1[5:0] ? myHhdoutVec_63 : _GEN_3783; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_20_T_1 = 16'h2b + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3786 = 6'h1 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3787 = 6'h2 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_2 : _GEN_3786; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3788 = 6'h3 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_3 : _GEN_3787; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3789 = 6'h4 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_4 : _GEN_3788; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3790 = 6'h5 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_5 : _GEN_3789; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3791 = 6'h6 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_6 : _GEN_3790; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3792 = 6'h7 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_7 : _GEN_3791; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3793 = 6'h8 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_8 : _GEN_3792; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3794 = 6'h9 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_9 : _GEN_3793; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3795 = 6'ha == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_10 : _GEN_3794; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3796 = 6'hb == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_11 : _GEN_3795; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3797 = 6'hc == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_12 : _GEN_3796; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3798 = 6'hd == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_13 : _GEN_3797; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3799 = 6'he == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_14 : _GEN_3798; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3800 = 6'hf == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_15 : _GEN_3799; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3801 = 6'h10 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_16 : _GEN_3800; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3802 = 6'h11 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_17 : _GEN_3801; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3803 = 6'h12 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_18 : _GEN_3802; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3804 = 6'h13 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_19 : _GEN_3803; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3805 = 6'h14 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_20 : _GEN_3804; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3806 = 6'h15 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_21 : _GEN_3805; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3807 = 6'h16 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_22 : _GEN_3806; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3808 = 6'h17 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_23 : _GEN_3807; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3809 = 6'h18 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_24 : _GEN_3808; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3810 = 6'h19 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_25 : _GEN_3809; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3811 = 6'h1a == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_26 : _GEN_3810; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3812 = 6'h1b == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_27 : _GEN_3811; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3813 = 6'h1c == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_28 : _GEN_3812; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3814 = 6'h1d == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_29 : _GEN_3813; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3815 = 6'h1e == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_30 : _GEN_3814; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3816 = 6'h1f == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_31 : _GEN_3815; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3817 = 6'h20 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_32 : _GEN_3816; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3818 = 6'h21 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_33 : _GEN_3817; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3819 = 6'h22 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_34 : _GEN_3818; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3820 = 6'h23 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_35 : _GEN_3819; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3821 = 6'h24 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_36 : _GEN_3820; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3822 = 6'h25 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_37 : _GEN_3821; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3823 = 6'h26 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_38 : _GEN_3822; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3824 = 6'h27 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_39 : _GEN_3823; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3825 = 6'h28 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_40 : _GEN_3824; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3826 = 6'h29 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_41 : _GEN_3825; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3827 = 6'h2a == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_42 : _GEN_3826; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3828 = 6'h2b == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_43 : _GEN_3827; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3829 = 6'h2c == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_44 : _GEN_3828; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3830 = 6'h2d == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_45 : _GEN_3829; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3831 = 6'h2e == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_46 : _GEN_3830; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3832 = 6'h2f == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_47 : _GEN_3831; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3833 = 6'h30 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_48 : _GEN_3832; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3834 = 6'h31 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_49 : _GEN_3833; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3835 = 6'h32 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_50 : _GEN_3834; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3836 = 6'h33 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_51 : _GEN_3835; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3837 = 6'h34 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_52 : _GEN_3836; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3838 = 6'h35 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_53 : _GEN_3837; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3839 = 6'h36 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_54 : _GEN_3838; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3840 = 6'h37 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_55 : _GEN_3839; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3841 = 6'h38 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_56 : _GEN_3840; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3842 = 6'h39 == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_57 : _GEN_3841; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3843 = 6'h3a == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_58 : _GEN_3842; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3844 = 6'h3b == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_59 : _GEN_3843; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3845 = 6'h3c == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_60 : _GEN_3844; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3846 = 6'h3d == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_61 : _GEN_3845; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3847 = 6'h3e == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_62 : _GEN_3846; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_20 = 6'h3f == _myHhdoutVec2_20_T_1[5:0] ? myHhdoutVec_63 : _GEN_3847; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_19_T_1 = 16'h2c + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3850 = 6'h1 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3851 = 6'h2 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_2 : _GEN_3850; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3852 = 6'h3 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_3 : _GEN_3851; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3853 = 6'h4 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_4 : _GEN_3852; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3854 = 6'h5 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_5 : _GEN_3853; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3855 = 6'h6 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_6 : _GEN_3854; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3856 = 6'h7 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_7 : _GEN_3855; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3857 = 6'h8 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_8 : _GEN_3856; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3858 = 6'h9 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_9 : _GEN_3857; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3859 = 6'ha == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_10 : _GEN_3858; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3860 = 6'hb == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_11 : _GEN_3859; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3861 = 6'hc == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_12 : _GEN_3860; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3862 = 6'hd == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_13 : _GEN_3861; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3863 = 6'he == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_14 : _GEN_3862; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3864 = 6'hf == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_15 : _GEN_3863; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3865 = 6'h10 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_16 : _GEN_3864; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3866 = 6'h11 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_17 : _GEN_3865; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3867 = 6'h12 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_18 : _GEN_3866; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3868 = 6'h13 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_19 : _GEN_3867; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3869 = 6'h14 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_20 : _GEN_3868; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3870 = 6'h15 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_21 : _GEN_3869; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3871 = 6'h16 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_22 : _GEN_3870; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3872 = 6'h17 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_23 : _GEN_3871; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3873 = 6'h18 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_24 : _GEN_3872; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3874 = 6'h19 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_25 : _GEN_3873; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3875 = 6'h1a == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_26 : _GEN_3874; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3876 = 6'h1b == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_27 : _GEN_3875; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3877 = 6'h1c == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_28 : _GEN_3876; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3878 = 6'h1d == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_29 : _GEN_3877; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3879 = 6'h1e == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_30 : _GEN_3878; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3880 = 6'h1f == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_31 : _GEN_3879; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3881 = 6'h20 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_32 : _GEN_3880; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3882 = 6'h21 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_33 : _GEN_3881; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3883 = 6'h22 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_34 : _GEN_3882; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3884 = 6'h23 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_35 : _GEN_3883; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3885 = 6'h24 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_36 : _GEN_3884; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3886 = 6'h25 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_37 : _GEN_3885; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3887 = 6'h26 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_38 : _GEN_3886; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3888 = 6'h27 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_39 : _GEN_3887; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3889 = 6'h28 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_40 : _GEN_3888; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3890 = 6'h29 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_41 : _GEN_3889; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3891 = 6'h2a == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_42 : _GEN_3890; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3892 = 6'h2b == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_43 : _GEN_3891; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3893 = 6'h2c == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_44 : _GEN_3892; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3894 = 6'h2d == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_45 : _GEN_3893; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3895 = 6'h2e == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_46 : _GEN_3894; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3896 = 6'h2f == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_47 : _GEN_3895; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3897 = 6'h30 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_48 : _GEN_3896; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3898 = 6'h31 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_49 : _GEN_3897; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3899 = 6'h32 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_50 : _GEN_3898; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3900 = 6'h33 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_51 : _GEN_3899; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3901 = 6'h34 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_52 : _GEN_3900; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3902 = 6'h35 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_53 : _GEN_3901; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3903 = 6'h36 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_54 : _GEN_3902; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3904 = 6'h37 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_55 : _GEN_3903; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3905 = 6'h38 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_56 : _GEN_3904; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3906 = 6'h39 == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_57 : _GEN_3905; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3907 = 6'h3a == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_58 : _GEN_3906; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3908 = 6'h3b == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_59 : _GEN_3907; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3909 = 6'h3c == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_60 : _GEN_3908; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3910 = 6'h3d == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_61 : _GEN_3909; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3911 = 6'h3e == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_62 : _GEN_3910; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_19 = 6'h3f == _myHhdoutVec2_19_T_1[5:0] ? myHhdoutVec_63 : _GEN_3911; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_18_T_1 = 16'h2d + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3914 = 6'h1 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3915 = 6'h2 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_2 : _GEN_3914; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3916 = 6'h3 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_3 : _GEN_3915; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3917 = 6'h4 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_4 : _GEN_3916; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3918 = 6'h5 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_5 : _GEN_3917; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3919 = 6'h6 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_6 : _GEN_3918; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3920 = 6'h7 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_7 : _GEN_3919; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3921 = 6'h8 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_8 : _GEN_3920; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3922 = 6'h9 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_9 : _GEN_3921; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3923 = 6'ha == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_10 : _GEN_3922; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3924 = 6'hb == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_11 : _GEN_3923; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3925 = 6'hc == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_12 : _GEN_3924; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3926 = 6'hd == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_13 : _GEN_3925; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3927 = 6'he == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_14 : _GEN_3926; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3928 = 6'hf == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_15 : _GEN_3927; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3929 = 6'h10 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_16 : _GEN_3928; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3930 = 6'h11 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_17 : _GEN_3929; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3931 = 6'h12 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_18 : _GEN_3930; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3932 = 6'h13 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_19 : _GEN_3931; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3933 = 6'h14 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_20 : _GEN_3932; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3934 = 6'h15 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_21 : _GEN_3933; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3935 = 6'h16 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_22 : _GEN_3934; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3936 = 6'h17 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_23 : _GEN_3935; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3937 = 6'h18 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_24 : _GEN_3936; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3938 = 6'h19 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_25 : _GEN_3937; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3939 = 6'h1a == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_26 : _GEN_3938; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3940 = 6'h1b == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_27 : _GEN_3939; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3941 = 6'h1c == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_28 : _GEN_3940; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3942 = 6'h1d == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_29 : _GEN_3941; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3943 = 6'h1e == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_30 : _GEN_3942; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3944 = 6'h1f == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_31 : _GEN_3943; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3945 = 6'h20 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_32 : _GEN_3944; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3946 = 6'h21 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_33 : _GEN_3945; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3947 = 6'h22 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_34 : _GEN_3946; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3948 = 6'h23 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_35 : _GEN_3947; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3949 = 6'h24 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_36 : _GEN_3948; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3950 = 6'h25 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_37 : _GEN_3949; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3951 = 6'h26 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_38 : _GEN_3950; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3952 = 6'h27 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_39 : _GEN_3951; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3953 = 6'h28 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_40 : _GEN_3952; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3954 = 6'h29 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_41 : _GEN_3953; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3955 = 6'h2a == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_42 : _GEN_3954; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3956 = 6'h2b == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_43 : _GEN_3955; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3957 = 6'h2c == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_44 : _GEN_3956; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3958 = 6'h2d == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_45 : _GEN_3957; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3959 = 6'h2e == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_46 : _GEN_3958; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3960 = 6'h2f == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_47 : _GEN_3959; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3961 = 6'h30 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_48 : _GEN_3960; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3962 = 6'h31 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_49 : _GEN_3961; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3963 = 6'h32 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_50 : _GEN_3962; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3964 = 6'h33 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_51 : _GEN_3963; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3965 = 6'h34 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_52 : _GEN_3964; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3966 = 6'h35 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_53 : _GEN_3965; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3967 = 6'h36 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_54 : _GEN_3966; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3968 = 6'h37 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_55 : _GEN_3967; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3969 = 6'h38 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_56 : _GEN_3968; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3970 = 6'h39 == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_57 : _GEN_3969; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3971 = 6'h3a == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_58 : _GEN_3970; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3972 = 6'h3b == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_59 : _GEN_3971; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3973 = 6'h3c == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_60 : _GEN_3972; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3974 = 6'h3d == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_61 : _GEN_3973; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3975 = 6'h3e == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_62 : _GEN_3974; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_18 = 6'h3f == _myHhdoutVec2_18_T_1[5:0] ? myHhdoutVec_63 : _GEN_3975; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_17_T_1 = 16'h2e + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_3978 = 6'h1 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3979 = 6'h2 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_2 : _GEN_3978; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3980 = 6'h3 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_3 : _GEN_3979; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3981 = 6'h4 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_4 : _GEN_3980; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3982 = 6'h5 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_5 : _GEN_3981; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3983 = 6'h6 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_6 : _GEN_3982; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3984 = 6'h7 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_7 : _GEN_3983; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3985 = 6'h8 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_8 : _GEN_3984; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3986 = 6'h9 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_9 : _GEN_3985; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3987 = 6'ha == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_10 : _GEN_3986; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3988 = 6'hb == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_11 : _GEN_3987; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3989 = 6'hc == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_12 : _GEN_3988; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3990 = 6'hd == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_13 : _GEN_3989; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3991 = 6'he == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_14 : _GEN_3990; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3992 = 6'hf == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_15 : _GEN_3991; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3993 = 6'h10 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_16 : _GEN_3992; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3994 = 6'h11 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_17 : _GEN_3993; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3995 = 6'h12 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_18 : _GEN_3994; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3996 = 6'h13 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_19 : _GEN_3995; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3997 = 6'h14 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_20 : _GEN_3996; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3998 = 6'h15 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_21 : _GEN_3997; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_3999 = 6'h16 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_22 : _GEN_3998; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4000 = 6'h17 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_23 : _GEN_3999; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4001 = 6'h18 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_24 : _GEN_4000; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4002 = 6'h19 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_25 : _GEN_4001; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4003 = 6'h1a == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_26 : _GEN_4002; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4004 = 6'h1b == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_27 : _GEN_4003; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4005 = 6'h1c == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_28 : _GEN_4004; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4006 = 6'h1d == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_29 : _GEN_4005; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4007 = 6'h1e == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_30 : _GEN_4006; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4008 = 6'h1f == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_31 : _GEN_4007; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4009 = 6'h20 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_32 : _GEN_4008; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4010 = 6'h21 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_33 : _GEN_4009; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4011 = 6'h22 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_34 : _GEN_4010; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4012 = 6'h23 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_35 : _GEN_4011; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4013 = 6'h24 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_36 : _GEN_4012; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4014 = 6'h25 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_37 : _GEN_4013; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4015 = 6'h26 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_38 : _GEN_4014; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4016 = 6'h27 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_39 : _GEN_4015; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4017 = 6'h28 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_40 : _GEN_4016; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4018 = 6'h29 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_41 : _GEN_4017; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4019 = 6'h2a == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_42 : _GEN_4018; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4020 = 6'h2b == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_43 : _GEN_4019; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4021 = 6'h2c == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_44 : _GEN_4020; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4022 = 6'h2d == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_45 : _GEN_4021; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4023 = 6'h2e == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_46 : _GEN_4022; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4024 = 6'h2f == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_47 : _GEN_4023; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4025 = 6'h30 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_48 : _GEN_4024; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4026 = 6'h31 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_49 : _GEN_4025; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4027 = 6'h32 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_50 : _GEN_4026; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4028 = 6'h33 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_51 : _GEN_4027; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4029 = 6'h34 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_52 : _GEN_4028; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4030 = 6'h35 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_53 : _GEN_4029; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4031 = 6'h36 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_54 : _GEN_4030; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4032 = 6'h37 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_55 : _GEN_4031; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4033 = 6'h38 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_56 : _GEN_4032; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4034 = 6'h39 == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_57 : _GEN_4033; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4035 = 6'h3a == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_58 : _GEN_4034; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4036 = 6'h3b == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_59 : _GEN_4035; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4037 = 6'h3c == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_60 : _GEN_4036; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4038 = 6'h3d == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_61 : _GEN_4037; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4039 = 6'h3e == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_62 : _GEN_4038; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_17 = 6'h3f == _myHhdoutVec2_17_T_1[5:0] ? myHhdoutVec_63 : _GEN_4039; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_16_T_1 = 16'h2f + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4042 = 6'h1 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4043 = 6'h2 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_2 : _GEN_4042; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4044 = 6'h3 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_3 : _GEN_4043; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4045 = 6'h4 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_4 : _GEN_4044; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4046 = 6'h5 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_5 : _GEN_4045; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4047 = 6'h6 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_6 : _GEN_4046; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4048 = 6'h7 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_7 : _GEN_4047; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4049 = 6'h8 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_8 : _GEN_4048; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4050 = 6'h9 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_9 : _GEN_4049; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4051 = 6'ha == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_10 : _GEN_4050; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4052 = 6'hb == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_11 : _GEN_4051; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4053 = 6'hc == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_12 : _GEN_4052; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4054 = 6'hd == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_13 : _GEN_4053; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4055 = 6'he == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_14 : _GEN_4054; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4056 = 6'hf == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_15 : _GEN_4055; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4057 = 6'h10 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_16 : _GEN_4056; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4058 = 6'h11 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_17 : _GEN_4057; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4059 = 6'h12 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_18 : _GEN_4058; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4060 = 6'h13 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_19 : _GEN_4059; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4061 = 6'h14 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_20 : _GEN_4060; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4062 = 6'h15 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_21 : _GEN_4061; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4063 = 6'h16 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_22 : _GEN_4062; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4064 = 6'h17 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_23 : _GEN_4063; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4065 = 6'h18 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_24 : _GEN_4064; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4066 = 6'h19 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_25 : _GEN_4065; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4067 = 6'h1a == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_26 : _GEN_4066; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4068 = 6'h1b == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_27 : _GEN_4067; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4069 = 6'h1c == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_28 : _GEN_4068; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4070 = 6'h1d == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_29 : _GEN_4069; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4071 = 6'h1e == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_30 : _GEN_4070; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4072 = 6'h1f == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_31 : _GEN_4071; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4073 = 6'h20 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_32 : _GEN_4072; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4074 = 6'h21 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_33 : _GEN_4073; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4075 = 6'h22 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_34 : _GEN_4074; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4076 = 6'h23 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_35 : _GEN_4075; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4077 = 6'h24 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_36 : _GEN_4076; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4078 = 6'h25 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_37 : _GEN_4077; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4079 = 6'h26 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_38 : _GEN_4078; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4080 = 6'h27 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_39 : _GEN_4079; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4081 = 6'h28 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_40 : _GEN_4080; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4082 = 6'h29 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_41 : _GEN_4081; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4083 = 6'h2a == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_42 : _GEN_4082; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4084 = 6'h2b == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_43 : _GEN_4083; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4085 = 6'h2c == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_44 : _GEN_4084; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4086 = 6'h2d == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_45 : _GEN_4085; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4087 = 6'h2e == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_46 : _GEN_4086; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4088 = 6'h2f == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_47 : _GEN_4087; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4089 = 6'h30 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_48 : _GEN_4088; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4090 = 6'h31 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_49 : _GEN_4089; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4091 = 6'h32 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_50 : _GEN_4090; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4092 = 6'h33 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_51 : _GEN_4091; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4093 = 6'h34 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_52 : _GEN_4092; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4094 = 6'h35 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_53 : _GEN_4093; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4095 = 6'h36 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_54 : _GEN_4094; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4096 = 6'h37 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_55 : _GEN_4095; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4097 = 6'h38 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_56 : _GEN_4096; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4098 = 6'h39 == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_57 : _GEN_4097; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4099 = 6'h3a == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_58 : _GEN_4098; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4100 = 6'h3b == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_59 : _GEN_4099; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4101 = 6'h3c == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_60 : _GEN_4100; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4102 = 6'h3d == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_61 : _GEN_4101; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4103 = 6'h3e == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_62 : _GEN_4102; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_16 = 6'h3f == _myHhdoutVec2_16_T_1[5:0] ? myHhdoutVec_63 : _GEN_4103; // @[hh_core.scala 149:{52,52}]
  wire [255:0] myHhdoutWire_lo_hi_lo = {myHhdoutVec2_23,myHhdoutVec2_22,myHhdoutVec2_21,myHhdoutVec2_20,myHhdoutVec2_19,
    myHhdoutVec2_18,myHhdoutVec2_17,myHhdoutVec2_16}; // @[hh_core.scala 153:42]
  wire [15:0] _myHhdoutVec2_15_T_1 = 16'h30 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4106 = 6'h1 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4107 = 6'h2 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_2 : _GEN_4106; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4108 = 6'h3 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_3 : _GEN_4107; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4109 = 6'h4 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_4 : _GEN_4108; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4110 = 6'h5 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_5 : _GEN_4109; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4111 = 6'h6 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_6 : _GEN_4110; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4112 = 6'h7 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_7 : _GEN_4111; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4113 = 6'h8 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_8 : _GEN_4112; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4114 = 6'h9 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_9 : _GEN_4113; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4115 = 6'ha == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_10 : _GEN_4114; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4116 = 6'hb == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_11 : _GEN_4115; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4117 = 6'hc == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_12 : _GEN_4116; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4118 = 6'hd == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_13 : _GEN_4117; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4119 = 6'he == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_14 : _GEN_4118; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4120 = 6'hf == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_15 : _GEN_4119; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4121 = 6'h10 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_16 : _GEN_4120; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4122 = 6'h11 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_17 : _GEN_4121; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4123 = 6'h12 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_18 : _GEN_4122; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4124 = 6'h13 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_19 : _GEN_4123; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4125 = 6'h14 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_20 : _GEN_4124; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4126 = 6'h15 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_21 : _GEN_4125; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4127 = 6'h16 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_22 : _GEN_4126; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4128 = 6'h17 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_23 : _GEN_4127; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4129 = 6'h18 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_24 : _GEN_4128; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4130 = 6'h19 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_25 : _GEN_4129; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4131 = 6'h1a == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_26 : _GEN_4130; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4132 = 6'h1b == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_27 : _GEN_4131; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4133 = 6'h1c == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_28 : _GEN_4132; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4134 = 6'h1d == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_29 : _GEN_4133; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4135 = 6'h1e == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_30 : _GEN_4134; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4136 = 6'h1f == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_31 : _GEN_4135; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4137 = 6'h20 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_32 : _GEN_4136; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4138 = 6'h21 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_33 : _GEN_4137; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4139 = 6'h22 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_34 : _GEN_4138; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4140 = 6'h23 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_35 : _GEN_4139; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4141 = 6'h24 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_36 : _GEN_4140; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4142 = 6'h25 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_37 : _GEN_4141; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4143 = 6'h26 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_38 : _GEN_4142; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4144 = 6'h27 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_39 : _GEN_4143; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4145 = 6'h28 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_40 : _GEN_4144; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4146 = 6'h29 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_41 : _GEN_4145; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4147 = 6'h2a == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_42 : _GEN_4146; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4148 = 6'h2b == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_43 : _GEN_4147; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4149 = 6'h2c == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_44 : _GEN_4148; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4150 = 6'h2d == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_45 : _GEN_4149; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4151 = 6'h2e == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_46 : _GEN_4150; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4152 = 6'h2f == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_47 : _GEN_4151; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4153 = 6'h30 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_48 : _GEN_4152; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4154 = 6'h31 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_49 : _GEN_4153; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4155 = 6'h32 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_50 : _GEN_4154; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4156 = 6'h33 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_51 : _GEN_4155; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4157 = 6'h34 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_52 : _GEN_4156; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4158 = 6'h35 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_53 : _GEN_4157; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4159 = 6'h36 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_54 : _GEN_4158; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4160 = 6'h37 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_55 : _GEN_4159; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4161 = 6'h38 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_56 : _GEN_4160; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4162 = 6'h39 == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_57 : _GEN_4161; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4163 = 6'h3a == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_58 : _GEN_4162; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4164 = 6'h3b == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_59 : _GEN_4163; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4165 = 6'h3c == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_60 : _GEN_4164; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4166 = 6'h3d == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_61 : _GEN_4165; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4167 = 6'h3e == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_62 : _GEN_4166; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_15 = 6'h3f == _myHhdoutVec2_15_T_1[5:0] ? myHhdoutVec_63 : _GEN_4167; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_14_T_1 = 16'h31 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4170 = 6'h1 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4171 = 6'h2 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_2 : _GEN_4170; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4172 = 6'h3 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_3 : _GEN_4171; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4173 = 6'h4 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_4 : _GEN_4172; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4174 = 6'h5 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_5 : _GEN_4173; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4175 = 6'h6 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_6 : _GEN_4174; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4176 = 6'h7 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_7 : _GEN_4175; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4177 = 6'h8 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_8 : _GEN_4176; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4178 = 6'h9 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_9 : _GEN_4177; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4179 = 6'ha == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_10 : _GEN_4178; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4180 = 6'hb == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_11 : _GEN_4179; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4181 = 6'hc == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_12 : _GEN_4180; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4182 = 6'hd == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_13 : _GEN_4181; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4183 = 6'he == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_14 : _GEN_4182; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4184 = 6'hf == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_15 : _GEN_4183; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4185 = 6'h10 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_16 : _GEN_4184; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4186 = 6'h11 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_17 : _GEN_4185; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4187 = 6'h12 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_18 : _GEN_4186; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4188 = 6'h13 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_19 : _GEN_4187; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4189 = 6'h14 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_20 : _GEN_4188; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4190 = 6'h15 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_21 : _GEN_4189; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4191 = 6'h16 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_22 : _GEN_4190; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4192 = 6'h17 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_23 : _GEN_4191; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4193 = 6'h18 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_24 : _GEN_4192; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4194 = 6'h19 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_25 : _GEN_4193; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4195 = 6'h1a == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_26 : _GEN_4194; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4196 = 6'h1b == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_27 : _GEN_4195; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4197 = 6'h1c == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_28 : _GEN_4196; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4198 = 6'h1d == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_29 : _GEN_4197; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4199 = 6'h1e == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_30 : _GEN_4198; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4200 = 6'h1f == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_31 : _GEN_4199; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4201 = 6'h20 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_32 : _GEN_4200; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4202 = 6'h21 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_33 : _GEN_4201; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4203 = 6'h22 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_34 : _GEN_4202; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4204 = 6'h23 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_35 : _GEN_4203; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4205 = 6'h24 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_36 : _GEN_4204; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4206 = 6'h25 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_37 : _GEN_4205; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4207 = 6'h26 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_38 : _GEN_4206; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4208 = 6'h27 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_39 : _GEN_4207; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4209 = 6'h28 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_40 : _GEN_4208; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4210 = 6'h29 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_41 : _GEN_4209; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4211 = 6'h2a == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_42 : _GEN_4210; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4212 = 6'h2b == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_43 : _GEN_4211; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4213 = 6'h2c == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_44 : _GEN_4212; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4214 = 6'h2d == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_45 : _GEN_4213; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4215 = 6'h2e == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_46 : _GEN_4214; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4216 = 6'h2f == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_47 : _GEN_4215; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4217 = 6'h30 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_48 : _GEN_4216; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4218 = 6'h31 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_49 : _GEN_4217; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4219 = 6'h32 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_50 : _GEN_4218; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4220 = 6'h33 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_51 : _GEN_4219; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4221 = 6'h34 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_52 : _GEN_4220; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4222 = 6'h35 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_53 : _GEN_4221; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4223 = 6'h36 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_54 : _GEN_4222; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4224 = 6'h37 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_55 : _GEN_4223; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4225 = 6'h38 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_56 : _GEN_4224; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4226 = 6'h39 == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_57 : _GEN_4225; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4227 = 6'h3a == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_58 : _GEN_4226; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4228 = 6'h3b == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_59 : _GEN_4227; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4229 = 6'h3c == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_60 : _GEN_4228; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4230 = 6'h3d == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_61 : _GEN_4229; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4231 = 6'h3e == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_62 : _GEN_4230; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_14 = 6'h3f == _myHhdoutVec2_14_T_1[5:0] ? myHhdoutVec_63 : _GEN_4231; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_13_T_1 = 16'h32 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4234 = 6'h1 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4235 = 6'h2 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_2 : _GEN_4234; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4236 = 6'h3 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_3 : _GEN_4235; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4237 = 6'h4 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_4 : _GEN_4236; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4238 = 6'h5 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_5 : _GEN_4237; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4239 = 6'h6 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_6 : _GEN_4238; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4240 = 6'h7 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_7 : _GEN_4239; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4241 = 6'h8 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_8 : _GEN_4240; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4242 = 6'h9 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_9 : _GEN_4241; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4243 = 6'ha == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_10 : _GEN_4242; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4244 = 6'hb == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_11 : _GEN_4243; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4245 = 6'hc == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_12 : _GEN_4244; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4246 = 6'hd == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_13 : _GEN_4245; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4247 = 6'he == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_14 : _GEN_4246; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4248 = 6'hf == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_15 : _GEN_4247; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4249 = 6'h10 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_16 : _GEN_4248; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4250 = 6'h11 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_17 : _GEN_4249; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4251 = 6'h12 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_18 : _GEN_4250; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4252 = 6'h13 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_19 : _GEN_4251; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4253 = 6'h14 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_20 : _GEN_4252; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4254 = 6'h15 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_21 : _GEN_4253; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4255 = 6'h16 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_22 : _GEN_4254; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4256 = 6'h17 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_23 : _GEN_4255; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4257 = 6'h18 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_24 : _GEN_4256; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4258 = 6'h19 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_25 : _GEN_4257; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4259 = 6'h1a == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_26 : _GEN_4258; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4260 = 6'h1b == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_27 : _GEN_4259; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4261 = 6'h1c == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_28 : _GEN_4260; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4262 = 6'h1d == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_29 : _GEN_4261; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4263 = 6'h1e == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_30 : _GEN_4262; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4264 = 6'h1f == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_31 : _GEN_4263; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4265 = 6'h20 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_32 : _GEN_4264; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4266 = 6'h21 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_33 : _GEN_4265; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4267 = 6'h22 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_34 : _GEN_4266; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4268 = 6'h23 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_35 : _GEN_4267; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4269 = 6'h24 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_36 : _GEN_4268; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4270 = 6'h25 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_37 : _GEN_4269; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4271 = 6'h26 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_38 : _GEN_4270; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4272 = 6'h27 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_39 : _GEN_4271; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4273 = 6'h28 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_40 : _GEN_4272; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4274 = 6'h29 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_41 : _GEN_4273; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4275 = 6'h2a == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_42 : _GEN_4274; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4276 = 6'h2b == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_43 : _GEN_4275; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4277 = 6'h2c == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_44 : _GEN_4276; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4278 = 6'h2d == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_45 : _GEN_4277; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4279 = 6'h2e == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_46 : _GEN_4278; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4280 = 6'h2f == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_47 : _GEN_4279; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4281 = 6'h30 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_48 : _GEN_4280; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4282 = 6'h31 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_49 : _GEN_4281; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4283 = 6'h32 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_50 : _GEN_4282; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4284 = 6'h33 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_51 : _GEN_4283; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4285 = 6'h34 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_52 : _GEN_4284; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4286 = 6'h35 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_53 : _GEN_4285; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4287 = 6'h36 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_54 : _GEN_4286; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4288 = 6'h37 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_55 : _GEN_4287; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4289 = 6'h38 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_56 : _GEN_4288; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4290 = 6'h39 == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_57 : _GEN_4289; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4291 = 6'h3a == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_58 : _GEN_4290; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4292 = 6'h3b == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_59 : _GEN_4291; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4293 = 6'h3c == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_60 : _GEN_4292; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4294 = 6'h3d == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_61 : _GEN_4293; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4295 = 6'h3e == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_62 : _GEN_4294; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_13 = 6'h3f == _myHhdoutVec2_13_T_1[5:0] ? myHhdoutVec_63 : _GEN_4295; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_12_T_1 = 16'h33 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4298 = 6'h1 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4299 = 6'h2 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_2 : _GEN_4298; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4300 = 6'h3 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_3 : _GEN_4299; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4301 = 6'h4 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_4 : _GEN_4300; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4302 = 6'h5 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_5 : _GEN_4301; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4303 = 6'h6 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_6 : _GEN_4302; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4304 = 6'h7 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_7 : _GEN_4303; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4305 = 6'h8 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_8 : _GEN_4304; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4306 = 6'h9 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_9 : _GEN_4305; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4307 = 6'ha == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_10 : _GEN_4306; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4308 = 6'hb == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_11 : _GEN_4307; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4309 = 6'hc == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_12 : _GEN_4308; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4310 = 6'hd == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_13 : _GEN_4309; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4311 = 6'he == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_14 : _GEN_4310; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4312 = 6'hf == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_15 : _GEN_4311; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4313 = 6'h10 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_16 : _GEN_4312; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4314 = 6'h11 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_17 : _GEN_4313; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4315 = 6'h12 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_18 : _GEN_4314; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4316 = 6'h13 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_19 : _GEN_4315; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4317 = 6'h14 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_20 : _GEN_4316; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4318 = 6'h15 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_21 : _GEN_4317; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4319 = 6'h16 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_22 : _GEN_4318; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4320 = 6'h17 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_23 : _GEN_4319; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4321 = 6'h18 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_24 : _GEN_4320; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4322 = 6'h19 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_25 : _GEN_4321; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4323 = 6'h1a == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_26 : _GEN_4322; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4324 = 6'h1b == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_27 : _GEN_4323; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4325 = 6'h1c == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_28 : _GEN_4324; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4326 = 6'h1d == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_29 : _GEN_4325; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4327 = 6'h1e == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_30 : _GEN_4326; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4328 = 6'h1f == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_31 : _GEN_4327; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4329 = 6'h20 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_32 : _GEN_4328; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4330 = 6'h21 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_33 : _GEN_4329; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4331 = 6'h22 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_34 : _GEN_4330; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4332 = 6'h23 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_35 : _GEN_4331; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4333 = 6'h24 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_36 : _GEN_4332; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4334 = 6'h25 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_37 : _GEN_4333; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4335 = 6'h26 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_38 : _GEN_4334; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4336 = 6'h27 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_39 : _GEN_4335; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4337 = 6'h28 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_40 : _GEN_4336; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4338 = 6'h29 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_41 : _GEN_4337; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4339 = 6'h2a == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_42 : _GEN_4338; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4340 = 6'h2b == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_43 : _GEN_4339; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4341 = 6'h2c == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_44 : _GEN_4340; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4342 = 6'h2d == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_45 : _GEN_4341; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4343 = 6'h2e == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_46 : _GEN_4342; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4344 = 6'h2f == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_47 : _GEN_4343; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4345 = 6'h30 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_48 : _GEN_4344; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4346 = 6'h31 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_49 : _GEN_4345; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4347 = 6'h32 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_50 : _GEN_4346; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4348 = 6'h33 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_51 : _GEN_4347; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4349 = 6'h34 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_52 : _GEN_4348; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4350 = 6'h35 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_53 : _GEN_4349; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4351 = 6'h36 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_54 : _GEN_4350; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4352 = 6'h37 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_55 : _GEN_4351; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4353 = 6'h38 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_56 : _GEN_4352; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4354 = 6'h39 == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_57 : _GEN_4353; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4355 = 6'h3a == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_58 : _GEN_4354; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4356 = 6'h3b == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_59 : _GEN_4355; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4357 = 6'h3c == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_60 : _GEN_4356; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4358 = 6'h3d == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_61 : _GEN_4357; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4359 = 6'h3e == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_62 : _GEN_4358; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_12 = 6'h3f == _myHhdoutVec2_12_T_1[5:0] ? myHhdoutVec_63 : _GEN_4359; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_11_T_1 = 16'h34 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4362 = 6'h1 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4363 = 6'h2 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_2 : _GEN_4362; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4364 = 6'h3 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_3 : _GEN_4363; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4365 = 6'h4 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_4 : _GEN_4364; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4366 = 6'h5 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_5 : _GEN_4365; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4367 = 6'h6 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_6 : _GEN_4366; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4368 = 6'h7 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_7 : _GEN_4367; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4369 = 6'h8 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_8 : _GEN_4368; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4370 = 6'h9 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_9 : _GEN_4369; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4371 = 6'ha == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_10 : _GEN_4370; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4372 = 6'hb == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_11 : _GEN_4371; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4373 = 6'hc == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_12 : _GEN_4372; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4374 = 6'hd == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_13 : _GEN_4373; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4375 = 6'he == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_14 : _GEN_4374; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4376 = 6'hf == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_15 : _GEN_4375; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4377 = 6'h10 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_16 : _GEN_4376; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4378 = 6'h11 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_17 : _GEN_4377; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4379 = 6'h12 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_18 : _GEN_4378; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4380 = 6'h13 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_19 : _GEN_4379; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4381 = 6'h14 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_20 : _GEN_4380; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4382 = 6'h15 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_21 : _GEN_4381; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4383 = 6'h16 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_22 : _GEN_4382; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4384 = 6'h17 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_23 : _GEN_4383; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4385 = 6'h18 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_24 : _GEN_4384; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4386 = 6'h19 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_25 : _GEN_4385; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4387 = 6'h1a == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_26 : _GEN_4386; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4388 = 6'h1b == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_27 : _GEN_4387; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4389 = 6'h1c == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_28 : _GEN_4388; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4390 = 6'h1d == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_29 : _GEN_4389; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4391 = 6'h1e == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_30 : _GEN_4390; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4392 = 6'h1f == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_31 : _GEN_4391; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4393 = 6'h20 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_32 : _GEN_4392; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4394 = 6'h21 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_33 : _GEN_4393; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4395 = 6'h22 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_34 : _GEN_4394; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4396 = 6'h23 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_35 : _GEN_4395; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4397 = 6'h24 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_36 : _GEN_4396; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4398 = 6'h25 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_37 : _GEN_4397; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4399 = 6'h26 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_38 : _GEN_4398; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4400 = 6'h27 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_39 : _GEN_4399; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4401 = 6'h28 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_40 : _GEN_4400; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4402 = 6'h29 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_41 : _GEN_4401; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4403 = 6'h2a == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_42 : _GEN_4402; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4404 = 6'h2b == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_43 : _GEN_4403; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4405 = 6'h2c == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_44 : _GEN_4404; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4406 = 6'h2d == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_45 : _GEN_4405; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4407 = 6'h2e == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_46 : _GEN_4406; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4408 = 6'h2f == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_47 : _GEN_4407; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4409 = 6'h30 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_48 : _GEN_4408; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4410 = 6'h31 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_49 : _GEN_4409; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4411 = 6'h32 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_50 : _GEN_4410; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4412 = 6'h33 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_51 : _GEN_4411; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4413 = 6'h34 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_52 : _GEN_4412; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4414 = 6'h35 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_53 : _GEN_4413; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4415 = 6'h36 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_54 : _GEN_4414; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4416 = 6'h37 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_55 : _GEN_4415; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4417 = 6'h38 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_56 : _GEN_4416; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4418 = 6'h39 == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_57 : _GEN_4417; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4419 = 6'h3a == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_58 : _GEN_4418; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4420 = 6'h3b == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_59 : _GEN_4419; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4421 = 6'h3c == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_60 : _GEN_4420; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4422 = 6'h3d == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_61 : _GEN_4421; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4423 = 6'h3e == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_62 : _GEN_4422; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_11 = 6'h3f == _myHhdoutVec2_11_T_1[5:0] ? myHhdoutVec_63 : _GEN_4423; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_10_T_1 = 16'h35 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4426 = 6'h1 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4427 = 6'h2 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_2 : _GEN_4426; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4428 = 6'h3 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_3 : _GEN_4427; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4429 = 6'h4 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_4 : _GEN_4428; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4430 = 6'h5 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_5 : _GEN_4429; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4431 = 6'h6 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_6 : _GEN_4430; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4432 = 6'h7 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_7 : _GEN_4431; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4433 = 6'h8 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_8 : _GEN_4432; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4434 = 6'h9 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_9 : _GEN_4433; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4435 = 6'ha == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_10 : _GEN_4434; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4436 = 6'hb == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_11 : _GEN_4435; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4437 = 6'hc == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_12 : _GEN_4436; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4438 = 6'hd == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_13 : _GEN_4437; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4439 = 6'he == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_14 : _GEN_4438; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4440 = 6'hf == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_15 : _GEN_4439; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4441 = 6'h10 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_16 : _GEN_4440; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4442 = 6'h11 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_17 : _GEN_4441; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4443 = 6'h12 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_18 : _GEN_4442; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4444 = 6'h13 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_19 : _GEN_4443; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4445 = 6'h14 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_20 : _GEN_4444; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4446 = 6'h15 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_21 : _GEN_4445; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4447 = 6'h16 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_22 : _GEN_4446; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4448 = 6'h17 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_23 : _GEN_4447; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4449 = 6'h18 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_24 : _GEN_4448; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4450 = 6'h19 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_25 : _GEN_4449; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4451 = 6'h1a == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_26 : _GEN_4450; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4452 = 6'h1b == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_27 : _GEN_4451; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4453 = 6'h1c == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_28 : _GEN_4452; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4454 = 6'h1d == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_29 : _GEN_4453; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4455 = 6'h1e == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_30 : _GEN_4454; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4456 = 6'h1f == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_31 : _GEN_4455; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4457 = 6'h20 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_32 : _GEN_4456; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4458 = 6'h21 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_33 : _GEN_4457; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4459 = 6'h22 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_34 : _GEN_4458; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4460 = 6'h23 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_35 : _GEN_4459; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4461 = 6'h24 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_36 : _GEN_4460; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4462 = 6'h25 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_37 : _GEN_4461; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4463 = 6'h26 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_38 : _GEN_4462; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4464 = 6'h27 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_39 : _GEN_4463; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4465 = 6'h28 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_40 : _GEN_4464; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4466 = 6'h29 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_41 : _GEN_4465; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4467 = 6'h2a == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_42 : _GEN_4466; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4468 = 6'h2b == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_43 : _GEN_4467; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4469 = 6'h2c == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_44 : _GEN_4468; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4470 = 6'h2d == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_45 : _GEN_4469; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4471 = 6'h2e == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_46 : _GEN_4470; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4472 = 6'h2f == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_47 : _GEN_4471; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4473 = 6'h30 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_48 : _GEN_4472; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4474 = 6'h31 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_49 : _GEN_4473; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4475 = 6'h32 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_50 : _GEN_4474; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4476 = 6'h33 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_51 : _GEN_4475; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4477 = 6'h34 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_52 : _GEN_4476; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4478 = 6'h35 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_53 : _GEN_4477; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4479 = 6'h36 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_54 : _GEN_4478; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4480 = 6'h37 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_55 : _GEN_4479; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4481 = 6'h38 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_56 : _GEN_4480; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4482 = 6'h39 == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_57 : _GEN_4481; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4483 = 6'h3a == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_58 : _GEN_4482; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4484 = 6'h3b == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_59 : _GEN_4483; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4485 = 6'h3c == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_60 : _GEN_4484; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4486 = 6'h3d == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_61 : _GEN_4485; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4487 = 6'h3e == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_62 : _GEN_4486; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_10 = 6'h3f == _myHhdoutVec2_10_T_1[5:0] ? myHhdoutVec_63 : _GEN_4487; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_9_T_1 = 16'h36 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4490 = 6'h1 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4491 = 6'h2 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_2 : _GEN_4490; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4492 = 6'h3 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_3 : _GEN_4491; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4493 = 6'h4 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_4 : _GEN_4492; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4494 = 6'h5 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_5 : _GEN_4493; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4495 = 6'h6 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_6 : _GEN_4494; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4496 = 6'h7 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_7 : _GEN_4495; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4497 = 6'h8 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_8 : _GEN_4496; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4498 = 6'h9 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_9 : _GEN_4497; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4499 = 6'ha == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_10 : _GEN_4498; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4500 = 6'hb == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_11 : _GEN_4499; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4501 = 6'hc == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_12 : _GEN_4500; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4502 = 6'hd == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_13 : _GEN_4501; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4503 = 6'he == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_14 : _GEN_4502; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4504 = 6'hf == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_15 : _GEN_4503; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4505 = 6'h10 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_16 : _GEN_4504; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4506 = 6'h11 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_17 : _GEN_4505; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4507 = 6'h12 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_18 : _GEN_4506; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4508 = 6'h13 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_19 : _GEN_4507; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4509 = 6'h14 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_20 : _GEN_4508; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4510 = 6'h15 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_21 : _GEN_4509; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4511 = 6'h16 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_22 : _GEN_4510; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4512 = 6'h17 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_23 : _GEN_4511; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4513 = 6'h18 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_24 : _GEN_4512; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4514 = 6'h19 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_25 : _GEN_4513; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4515 = 6'h1a == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_26 : _GEN_4514; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4516 = 6'h1b == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_27 : _GEN_4515; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4517 = 6'h1c == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_28 : _GEN_4516; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4518 = 6'h1d == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_29 : _GEN_4517; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4519 = 6'h1e == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_30 : _GEN_4518; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4520 = 6'h1f == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_31 : _GEN_4519; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4521 = 6'h20 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_32 : _GEN_4520; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4522 = 6'h21 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_33 : _GEN_4521; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4523 = 6'h22 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_34 : _GEN_4522; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4524 = 6'h23 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_35 : _GEN_4523; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4525 = 6'h24 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_36 : _GEN_4524; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4526 = 6'h25 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_37 : _GEN_4525; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4527 = 6'h26 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_38 : _GEN_4526; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4528 = 6'h27 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_39 : _GEN_4527; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4529 = 6'h28 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_40 : _GEN_4528; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4530 = 6'h29 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_41 : _GEN_4529; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4531 = 6'h2a == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_42 : _GEN_4530; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4532 = 6'h2b == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_43 : _GEN_4531; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4533 = 6'h2c == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_44 : _GEN_4532; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4534 = 6'h2d == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_45 : _GEN_4533; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4535 = 6'h2e == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_46 : _GEN_4534; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4536 = 6'h2f == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_47 : _GEN_4535; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4537 = 6'h30 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_48 : _GEN_4536; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4538 = 6'h31 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_49 : _GEN_4537; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4539 = 6'h32 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_50 : _GEN_4538; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4540 = 6'h33 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_51 : _GEN_4539; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4541 = 6'h34 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_52 : _GEN_4540; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4542 = 6'h35 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_53 : _GEN_4541; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4543 = 6'h36 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_54 : _GEN_4542; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4544 = 6'h37 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_55 : _GEN_4543; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4545 = 6'h38 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_56 : _GEN_4544; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4546 = 6'h39 == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_57 : _GEN_4545; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4547 = 6'h3a == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_58 : _GEN_4546; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4548 = 6'h3b == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_59 : _GEN_4547; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4549 = 6'h3c == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_60 : _GEN_4548; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4550 = 6'h3d == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_61 : _GEN_4549; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4551 = 6'h3e == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_62 : _GEN_4550; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_9 = 6'h3f == _myHhdoutVec2_9_T_1[5:0] ? myHhdoutVec_63 : _GEN_4551; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_8_T_1 = 16'h37 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4554 = 6'h1 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4555 = 6'h2 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_2 : _GEN_4554; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4556 = 6'h3 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_3 : _GEN_4555; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4557 = 6'h4 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_4 : _GEN_4556; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4558 = 6'h5 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_5 : _GEN_4557; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4559 = 6'h6 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_6 : _GEN_4558; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4560 = 6'h7 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_7 : _GEN_4559; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4561 = 6'h8 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_8 : _GEN_4560; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4562 = 6'h9 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_9 : _GEN_4561; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4563 = 6'ha == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_10 : _GEN_4562; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4564 = 6'hb == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_11 : _GEN_4563; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4565 = 6'hc == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_12 : _GEN_4564; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4566 = 6'hd == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_13 : _GEN_4565; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4567 = 6'he == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_14 : _GEN_4566; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4568 = 6'hf == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_15 : _GEN_4567; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4569 = 6'h10 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_16 : _GEN_4568; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4570 = 6'h11 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_17 : _GEN_4569; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4571 = 6'h12 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_18 : _GEN_4570; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4572 = 6'h13 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_19 : _GEN_4571; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4573 = 6'h14 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_20 : _GEN_4572; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4574 = 6'h15 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_21 : _GEN_4573; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4575 = 6'h16 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_22 : _GEN_4574; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4576 = 6'h17 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_23 : _GEN_4575; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4577 = 6'h18 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_24 : _GEN_4576; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4578 = 6'h19 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_25 : _GEN_4577; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4579 = 6'h1a == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_26 : _GEN_4578; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4580 = 6'h1b == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_27 : _GEN_4579; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4581 = 6'h1c == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_28 : _GEN_4580; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4582 = 6'h1d == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_29 : _GEN_4581; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4583 = 6'h1e == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_30 : _GEN_4582; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4584 = 6'h1f == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_31 : _GEN_4583; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4585 = 6'h20 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_32 : _GEN_4584; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4586 = 6'h21 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_33 : _GEN_4585; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4587 = 6'h22 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_34 : _GEN_4586; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4588 = 6'h23 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_35 : _GEN_4587; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4589 = 6'h24 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_36 : _GEN_4588; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4590 = 6'h25 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_37 : _GEN_4589; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4591 = 6'h26 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_38 : _GEN_4590; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4592 = 6'h27 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_39 : _GEN_4591; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4593 = 6'h28 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_40 : _GEN_4592; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4594 = 6'h29 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_41 : _GEN_4593; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4595 = 6'h2a == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_42 : _GEN_4594; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4596 = 6'h2b == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_43 : _GEN_4595; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4597 = 6'h2c == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_44 : _GEN_4596; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4598 = 6'h2d == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_45 : _GEN_4597; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4599 = 6'h2e == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_46 : _GEN_4598; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4600 = 6'h2f == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_47 : _GEN_4599; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4601 = 6'h30 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_48 : _GEN_4600; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4602 = 6'h31 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_49 : _GEN_4601; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4603 = 6'h32 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_50 : _GEN_4602; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4604 = 6'h33 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_51 : _GEN_4603; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4605 = 6'h34 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_52 : _GEN_4604; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4606 = 6'h35 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_53 : _GEN_4605; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4607 = 6'h36 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_54 : _GEN_4606; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4608 = 6'h37 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_55 : _GEN_4607; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4609 = 6'h38 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_56 : _GEN_4608; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4610 = 6'h39 == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_57 : _GEN_4609; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4611 = 6'h3a == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_58 : _GEN_4610; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4612 = 6'h3b == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_59 : _GEN_4611; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4613 = 6'h3c == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_60 : _GEN_4612; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4614 = 6'h3d == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_61 : _GEN_4613; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4615 = 6'h3e == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_62 : _GEN_4614; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_8 = 6'h3f == _myHhdoutVec2_8_T_1[5:0] ? myHhdoutVec_63 : _GEN_4615; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_7_T_1 = 16'h38 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4618 = 6'h1 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4619 = 6'h2 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_2 : _GEN_4618; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4620 = 6'h3 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_3 : _GEN_4619; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4621 = 6'h4 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_4 : _GEN_4620; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4622 = 6'h5 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_5 : _GEN_4621; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4623 = 6'h6 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_6 : _GEN_4622; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4624 = 6'h7 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_7 : _GEN_4623; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4625 = 6'h8 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_8 : _GEN_4624; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4626 = 6'h9 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_9 : _GEN_4625; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4627 = 6'ha == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_10 : _GEN_4626; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4628 = 6'hb == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_11 : _GEN_4627; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4629 = 6'hc == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_12 : _GEN_4628; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4630 = 6'hd == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_13 : _GEN_4629; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4631 = 6'he == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_14 : _GEN_4630; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4632 = 6'hf == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_15 : _GEN_4631; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4633 = 6'h10 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_16 : _GEN_4632; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4634 = 6'h11 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_17 : _GEN_4633; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4635 = 6'h12 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_18 : _GEN_4634; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4636 = 6'h13 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_19 : _GEN_4635; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4637 = 6'h14 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_20 : _GEN_4636; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4638 = 6'h15 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_21 : _GEN_4637; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4639 = 6'h16 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_22 : _GEN_4638; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4640 = 6'h17 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_23 : _GEN_4639; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4641 = 6'h18 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_24 : _GEN_4640; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4642 = 6'h19 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_25 : _GEN_4641; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4643 = 6'h1a == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_26 : _GEN_4642; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4644 = 6'h1b == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_27 : _GEN_4643; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4645 = 6'h1c == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_28 : _GEN_4644; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4646 = 6'h1d == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_29 : _GEN_4645; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4647 = 6'h1e == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_30 : _GEN_4646; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4648 = 6'h1f == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_31 : _GEN_4647; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4649 = 6'h20 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_32 : _GEN_4648; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4650 = 6'h21 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_33 : _GEN_4649; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4651 = 6'h22 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_34 : _GEN_4650; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4652 = 6'h23 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_35 : _GEN_4651; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4653 = 6'h24 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_36 : _GEN_4652; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4654 = 6'h25 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_37 : _GEN_4653; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4655 = 6'h26 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_38 : _GEN_4654; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4656 = 6'h27 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_39 : _GEN_4655; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4657 = 6'h28 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_40 : _GEN_4656; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4658 = 6'h29 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_41 : _GEN_4657; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4659 = 6'h2a == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_42 : _GEN_4658; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4660 = 6'h2b == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_43 : _GEN_4659; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4661 = 6'h2c == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_44 : _GEN_4660; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4662 = 6'h2d == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_45 : _GEN_4661; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4663 = 6'h2e == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_46 : _GEN_4662; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4664 = 6'h2f == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_47 : _GEN_4663; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4665 = 6'h30 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_48 : _GEN_4664; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4666 = 6'h31 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_49 : _GEN_4665; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4667 = 6'h32 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_50 : _GEN_4666; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4668 = 6'h33 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_51 : _GEN_4667; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4669 = 6'h34 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_52 : _GEN_4668; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4670 = 6'h35 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_53 : _GEN_4669; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4671 = 6'h36 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_54 : _GEN_4670; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4672 = 6'h37 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_55 : _GEN_4671; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4673 = 6'h38 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_56 : _GEN_4672; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4674 = 6'h39 == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_57 : _GEN_4673; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4675 = 6'h3a == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_58 : _GEN_4674; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4676 = 6'h3b == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_59 : _GEN_4675; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4677 = 6'h3c == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_60 : _GEN_4676; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4678 = 6'h3d == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_61 : _GEN_4677; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4679 = 6'h3e == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_62 : _GEN_4678; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_7 = 6'h3f == _myHhdoutVec2_7_T_1[5:0] ? myHhdoutVec_63 : _GEN_4679; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_6_T_1 = 16'h39 + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4682 = 6'h1 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4683 = 6'h2 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_2 : _GEN_4682; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4684 = 6'h3 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_3 : _GEN_4683; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4685 = 6'h4 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_4 : _GEN_4684; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4686 = 6'h5 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_5 : _GEN_4685; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4687 = 6'h6 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_6 : _GEN_4686; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4688 = 6'h7 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_7 : _GEN_4687; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4689 = 6'h8 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_8 : _GEN_4688; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4690 = 6'h9 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_9 : _GEN_4689; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4691 = 6'ha == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_10 : _GEN_4690; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4692 = 6'hb == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_11 : _GEN_4691; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4693 = 6'hc == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_12 : _GEN_4692; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4694 = 6'hd == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_13 : _GEN_4693; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4695 = 6'he == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_14 : _GEN_4694; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4696 = 6'hf == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_15 : _GEN_4695; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4697 = 6'h10 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_16 : _GEN_4696; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4698 = 6'h11 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_17 : _GEN_4697; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4699 = 6'h12 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_18 : _GEN_4698; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4700 = 6'h13 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_19 : _GEN_4699; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4701 = 6'h14 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_20 : _GEN_4700; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4702 = 6'h15 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_21 : _GEN_4701; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4703 = 6'h16 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_22 : _GEN_4702; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4704 = 6'h17 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_23 : _GEN_4703; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4705 = 6'h18 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_24 : _GEN_4704; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4706 = 6'h19 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_25 : _GEN_4705; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4707 = 6'h1a == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_26 : _GEN_4706; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4708 = 6'h1b == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_27 : _GEN_4707; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4709 = 6'h1c == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_28 : _GEN_4708; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4710 = 6'h1d == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_29 : _GEN_4709; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4711 = 6'h1e == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_30 : _GEN_4710; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4712 = 6'h1f == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_31 : _GEN_4711; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4713 = 6'h20 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_32 : _GEN_4712; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4714 = 6'h21 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_33 : _GEN_4713; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4715 = 6'h22 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_34 : _GEN_4714; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4716 = 6'h23 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_35 : _GEN_4715; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4717 = 6'h24 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_36 : _GEN_4716; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4718 = 6'h25 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_37 : _GEN_4717; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4719 = 6'h26 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_38 : _GEN_4718; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4720 = 6'h27 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_39 : _GEN_4719; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4721 = 6'h28 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_40 : _GEN_4720; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4722 = 6'h29 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_41 : _GEN_4721; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4723 = 6'h2a == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_42 : _GEN_4722; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4724 = 6'h2b == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_43 : _GEN_4723; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4725 = 6'h2c == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_44 : _GEN_4724; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4726 = 6'h2d == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_45 : _GEN_4725; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4727 = 6'h2e == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_46 : _GEN_4726; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4728 = 6'h2f == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_47 : _GEN_4727; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4729 = 6'h30 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_48 : _GEN_4728; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4730 = 6'h31 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_49 : _GEN_4729; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4731 = 6'h32 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_50 : _GEN_4730; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4732 = 6'h33 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_51 : _GEN_4731; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4733 = 6'h34 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_52 : _GEN_4732; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4734 = 6'h35 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_53 : _GEN_4733; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4735 = 6'h36 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_54 : _GEN_4734; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4736 = 6'h37 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_55 : _GEN_4735; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4737 = 6'h38 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_56 : _GEN_4736; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4738 = 6'h39 == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_57 : _GEN_4737; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4739 = 6'h3a == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_58 : _GEN_4738; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4740 = 6'h3b == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_59 : _GEN_4739; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4741 = 6'h3c == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_60 : _GEN_4740; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4742 = 6'h3d == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_61 : _GEN_4741; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4743 = 6'h3e == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_62 : _GEN_4742; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_6 = 6'h3f == _myHhdoutVec2_6_T_1[5:0] ? myHhdoutVec_63 : _GEN_4743; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_5_T_1 = 16'h3a + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4746 = 6'h1 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4747 = 6'h2 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_2 : _GEN_4746; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4748 = 6'h3 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_3 : _GEN_4747; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4749 = 6'h4 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_4 : _GEN_4748; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4750 = 6'h5 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_5 : _GEN_4749; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4751 = 6'h6 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_6 : _GEN_4750; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4752 = 6'h7 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_7 : _GEN_4751; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4753 = 6'h8 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_8 : _GEN_4752; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4754 = 6'h9 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_9 : _GEN_4753; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4755 = 6'ha == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_10 : _GEN_4754; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4756 = 6'hb == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_11 : _GEN_4755; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4757 = 6'hc == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_12 : _GEN_4756; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4758 = 6'hd == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_13 : _GEN_4757; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4759 = 6'he == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_14 : _GEN_4758; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4760 = 6'hf == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_15 : _GEN_4759; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4761 = 6'h10 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_16 : _GEN_4760; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4762 = 6'h11 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_17 : _GEN_4761; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4763 = 6'h12 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_18 : _GEN_4762; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4764 = 6'h13 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_19 : _GEN_4763; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4765 = 6'h14 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_20 : _GEN_4764; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4766 = 6'h15 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_21 : _GEN_4765; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4767 = 6'h16 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_22 : _GEN_4766; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4768 = 6'h17 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_23 : _GEN_4767; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4769 = 6'h18 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_24 : _GEN_4768; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4770 = 6'h19 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_25 : _GEN_4769; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4771 = 6'h1a == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_26 : _GEN_4770; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4772 = 6'h1b == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_27 : _GEN_4771; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4773 = 6'h1c == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_28 : _GEN_4772; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4774 = 6'h1d == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_29 : _GEN_4773; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4775 = 6'h1e == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_30 : _GEN_4774; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4776 = 6'h1f == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_31 : _GEN_4775; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4777 = 6'h20 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_32 : _GEN_4776; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4778 = 6'h21 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_33 : _GEN_4777; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4779 = 6'h22 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_34 : _GEN_4778; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4780 = 6'h23 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_35 : _GEN_4779; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4781 = 6'h24 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_36 : _GEN_4780; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4782 = 6'h25 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_37 : _GEN_4781; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4783 = 6'h26 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_38 : _GEN_4782; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4784 = 6'h27 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_39 : _GEN_4783; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4785 = 6'h28 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_40 : _GEN_4784; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4786 = 6'h29 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_41 : _GEN_4785; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4787 = 6'h2a == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_42 : _GEN_4786; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4788 = 6'h2b == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_43 : _GEN_4787; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4789 = 6'h2c == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_44 : _GEN_4788; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4790 = 6'h2d == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_45 : _GEN_4789; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4791 = 6'h2e == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_46 : _GEN_4790; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4792 = 6'h2f == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_47 : _GEN_4791; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4793 = 6'h30 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_48 : _GEN_4792; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4794 = 6'h31 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_49 : _GEN_4793; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4795 = 6'h32 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_50 : _GEN_4794; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4796 = 6'h33 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_51 : _GEN_4795; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4797 = 6'h34 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_52 : _GEN_4796; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4798 = 6'h35 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_53 : _GEN_4797; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4799 = 6'h36 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_54 : _GEN_4798; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4800 = 6'h37 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_55 : _GEN_4799; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4801 = 6'h38 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_56 : _GEN_4800; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4802 = 6'h39 == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_57 : _GEN_4801; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4803 = 6'h3a == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_58 : _GEN_4802; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4804 = 6'h3b == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_59 : _GEN_4803; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4805 = 6'h3c == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_60 : _GEN_4804; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4806 = 6'h3d == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_61 : _GEN_4805; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4807 = 6'h3e == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_62 : _GEN_4806; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_5 = 6'h3f == _myHhdoutVec2_5_T_1[5:0] ? myHhdoutVec_63 : _GEN_4807; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_4_T_1 = 16'h3b + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4810 = 6'h1 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4811 = 6'h2 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_2 : _GEN_4810; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4812 = 6'h3 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_3 : _GEN_4811; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4813 = 6'h4 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_4 : _GEN_4812; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4814 = 6'h5 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_5 : _GEN_4813; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4815 = 6'h6 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_6 : _GEN_4814; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4816 = 6'h7 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_7 : _GEN_4815; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4817 = 6'h8 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_8 : _GEN_4816; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4818 = 6'h9 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_9 : _GEN_4817; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4819 = 6'ha == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_10 : _GEN_4818; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4820 = 6'hb == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_11 : _GEN_4819; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4821 = 6'hc == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_12 : _GEN_4820; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4822 = 6'hd == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_13 : _GEN_4821; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4823 = 6'he == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_14 : _GEN_4822; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4824 = 6'hf == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_15 : _GEN_4823; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4825 = 6'h10 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_16 : _GEN_4824; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4826 = 6'h11 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_17 : _GEN_4825; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4827 = 6'h12 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_18 : _GEN_4826; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4828 = 6'h13 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_19 : _GEN_4827; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4829 = 6'h14 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_20 : _GEN_4828; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4830 = 6'h15 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_21 : _GEN_4829; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4831 = 6'h16 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_22 : _GEN_4830; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4832 = 6'h17 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_23 : _GEN_4831; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4833 = 6'h18 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_24 : _GEN_4832; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4834 = 6'h19 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_25 : _GEN_4833; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4835 = 6'h1a == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_26 : _GEN_4834; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4836 = 6'h1b == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_27 : _GEN_4835; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4837 = 6'h1c == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_28 : _GEN_4836; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4838 = 6'h1d == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_29 : _GEN_4837; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4839 = 6'h1e == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_30 : _GEN_4838; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4840 = 6'h1f == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_31 : _GEN_4839; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4841 = 6'h20 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_32 : _GEN_4840; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4842 = 6'h21 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_33 : _GEN_4841; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4843 = 6'h22 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_34 : _GEN_4842; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4844 = 6'h23 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_35 : _GEN_4843; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4845 = 6'h24 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_36 : _GEN_4844; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4846 = 6'h25 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_37 : _GEN_4845; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4847 = 6'h26 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_38 : _GEN_4846; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4848 = 6'h27 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_39 : _GEN_4847; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4849 = 6'h28 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_40 : _GEN_4848; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4850 = 6'h29 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_41 : _GEN_4849; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4851 = 6'h2a == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_42 : _GEN_4850; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4852 = 6'h2b == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_43 : _GEN_4851; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4853 = 6'h2c == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_44 : _GEN_4852; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4854 = 6'h2d == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_45 : _GEN_4853; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4855 = 6'h2e == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_46 : _GEN_4854; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4856 = 6'h2f == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_47 : _GEN_4855; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4857 = 6'h30 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_48 : _GEN_4856; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4858 = 6'h31 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_49 : _GEN_4857; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4859 = 6'h32 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_50 : _GEN_4858; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4860 = 6'h33 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_51 : _GEN_4859; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4861 = 6'h34 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_52 : _GEN_4860; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4862 = 6'h35 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_53 : _GEN_4861; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4863 = 6'h36 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_54 : _GEN_4862; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4864 = 6'h37 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_55 : _GEN_4863; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4865 = 6'h38 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_56 : _GEN_4864; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4866 = 6'h39 == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_57 : _GEN_4865; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4867 = 6'h3a == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_58 : _GEN_4866; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4868 = 6'h3b == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_59 : _GEN_4867; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4869 = 6'h3c == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_60 : _GEN_4868; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4870 = 6'h3d == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_61 : _GEN_4869; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4871 = 6'h3e == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_62 : _GEN_4870; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_4 = 6'h3f == _myHhdoutVec2_4_T_1[5:0] ? myHhdoutVec_63 : _GEN_4871; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_3_T_1 = 16'h3c + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4874 = 6'h1 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4875 = 6'h2 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_2 : _GEN_4874; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4876 = 6'h3 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_3 : _GEN_4875; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4877 = 6'h4 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_4 : _GEN_4876; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4878 = 6'h5 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_5 : _GEN_4877; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4879 = 6'h6 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_6 : _GEN_4878; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4880 = 6'h7 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_7 : _GEN_4879; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4881 = 6'h8 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_8 : _GEN_4880; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4882 = 6'h9 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_9 : _GEN_4881; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4883 = 6'ha == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_10 : _GEN_4882; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4884 = 6'hb == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_11 : _GEN_4883; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4885 = 6'hc == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_12 : _GEN_4884; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4886 = 6'hd == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_13 : _GEN_4885; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4887 = 6'he == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_14 : _GEN_4886; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4888 = 6'hf == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_15 : _GEN_4887; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4889 = 6'h10 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_16 : _GEN_4888; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4890 = 6'h11 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_17 : _GEN_4889; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4891 = 6'h12 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_18 : _GEN_4890; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4892 = 6'h13 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_19 : _GEN_4891; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4893 = 6'h14 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_20 : _GEN_4892; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4894 = 6'h15 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_21 : _GEN_4893; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4895 = 6'h16 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_22 : _GEN_4894; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4896 = 6'h17 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_23 : _GEN_4895; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4897 = 6'h18 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_24 : _GEN_4896; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4898 = 6'h19 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_25 : _GEN_4897; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4899 = 6'h1a == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_26 : _GEN_4898; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4900 = 6'h1b == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_27 : _GEN_4899; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4901 = 6'h1c == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_28 : _GEN_4900; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4902 = 6'h1d == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_29 : _GEN_4901; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4903 = 6'h1e == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_30 : _GEN_4902; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4904 = 6'h1f == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_31 : _GEN_4903; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4905 = 6'h20 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_32 : _GEN_4904; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4906 = 6'h21 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_33 : _GEN_4905; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4907 = 6'h22 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_34 : _GEN_4906; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4908 = 6'h23 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_35 : _GEN_4907; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4909 = 6'h24 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_36 : _GEN_4908; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4910 = 6'h25 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_37 : _GEN_4909; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4911 = 6'h26 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_38 : _GEN_4910; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4912 = 6'h27 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_39 : _GEN_4911; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4913 = 6'h28 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_40 : _GEN_4912; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4914 = 6'h29 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_41 : _GEN_4913; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4915 = 6'h2a == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_42 : _GEN_4914; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4916 = 6'h2b == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_43 : _GEN_4915; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4917 = 6'h2c == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_44 : _GEN_4916; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4918 = 6'h2d == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_45 : _GEN_4917; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4919 = 6'h2e == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_46 : _GEN_4918; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4920 = 6'h2f == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_47 : _GEN_4919; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4921 = 6'h30 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_48 : _GEN_4920; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4922 = 6'h31 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_49 : _GEN_4921; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4923 = 6'h32 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_50 : _GEN_4922; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4924 = 6'h33 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_51 : _GEN_4923; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4925 = 6'h34 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_52 : _GEN_4924; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4926 = 6'h35 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_53 : _GEN_4925; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4927 = 6'h36 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_54 : _GEN_4926; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4928 = 6'h37 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_55 : _GEN_4927; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4929 = 6'h38 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_56 : _GEN_4928; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4930 = 6'h39 == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_57 : _GEN_4929; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4931 = 6'h3a == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_58 : _GEN_4930; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4932 = 6'h3b == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_59 : _GEN_4931; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4933 = 6'h3c == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_60 : _GEN_4932; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4934 = 6'h3d == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_61 : _GEN_4933; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4935 = 6'h3e == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_62 : _GEN_4934; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_3 = 6'h3f == _myHhdoutVec2_3_T_1[5:0] ? myHhdoutVec_63 : _GEN_4935; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_2_T_1 = 16'h3d + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_4938 = 6'h1 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4939 = 6'h2 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_2 : _GEN_4938; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4940 = 6'h3 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_3 : _GEN_4939; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4941 = 6'h4 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_4 : _GEN_4940; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4942 = 6'h5 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_5 : _GEN_4941; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4943 = 6'h6 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_6 : _GEN_4942; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4944 = 6'h7 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_7 : _GEN_4943; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4945 = 6'h8 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_8 : _GEN_4944; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4946 = 6'h9 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_9 : _GEN_4945; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4947 = 6'ha == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_10 : _GEN_4946; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4948 = 6'hb == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_11 : _GEN_4947; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4949 = 6'hc == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_12 : _GEN_4948; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4950 = 6'hd == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_13 : _GEN_4949; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4951 = 6'he == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_14 : _GEN_4950; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4952 = 6'hf == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_15 : _GEN_4951; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4953 = 6'h10 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_16 : _GEN_4952; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4954 = 6'h11 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_17 : _GEN_4953; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4955 = 6'h12 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_18 : _GEN_4954; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4956 = 6'h13 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_19 : _GEN_4955; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4957 = 6'h14 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_20 : _GEN_4956; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4958 = 6'h15 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_21 : _GEN_4957; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4959 = 6'h16 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_22 : _GEN_4958; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4960 = 6'h17 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_23 : _GEN_4959; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4961 = 6'h18 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_24 : _GEN_4960; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4962 = 6'h19 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_25 : _GEN_4961; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4963 = 6'h1a == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_26 : _GEN_4962; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4964 = 6'h1b == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_27 : _GEN_4963; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4965 = 6'h1c == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_28 : _GEN_4964; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4966 = 6'h1d == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_29 : _GEN_4965; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4967 = 6'h1e == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_30 : _GEN_4966; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4968 = 6'h1f == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_31 : _GEN_4967; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4969 = 6'h20 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_32 : _GEN_4968; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4970 = 6'h21 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_33 : _GEN_4969; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4971 = 6'h22 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_34 : _GEN_4970; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4972 = 6'h23 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_35 : _GEN_4971; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4973 = 6'h24 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_36 : _GEN_4972; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4974 = 6'h25 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_37 : _GEN_4973; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4975 = 6'h26 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_38 : _GEN_4974; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4976 = 6'h27 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_39 : _GEN_4975; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4977 = 6'h28 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_40 : _GEN_4976; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4978 = 6'h29 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_41 : _GEN_4977; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4979 = 6'h2a == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_42 : _GEN_4978; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4980 = 6'h2b == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_43 : _GEN_4979; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4981 = 6'h2c == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_44 : _GEN_4980; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4982 = 6'h2d == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_45 : _GEN_4981; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4983 = 6'h2e == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_46 : _GEN_4982; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4984 = 6'h2f == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_47 : _GEN_4983; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4985 = 6'h30 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_48 : _GEN_4984; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4986 = 6'h31 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_49 : _GEN_4985; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4987 = 6'h32 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_50 : _GEN_4986; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4988 = 6'h33 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_51 : _GEN_4987; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4989 = 6'h34 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_52 : _GEN_4988; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4990 = 6'h35 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_53 : _GEN_4989; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4991 = 6'h36 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_54 : _GEN_4990; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4992 = 6'h37 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_55 : _GEN_4991; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4993 = 6'h38 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_56 : _GEN_4992; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4994 = 6'h39 == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_57 : _GEN_4993; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4995 = 6'h3a == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_58 : _GEN_4994; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4996 = 6'h3b == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_59 : _GEN_4995; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4997 = 6'h3c == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_60 : _GEN_4996; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4998 = 6'h3d == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_61 : _GEN_4997; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_4999 = 6'h3e == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_62 : _GEN_4998; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_2 = 6'h3f == _myHhdoutVec2_2_T_1[5:0] ? myHhdoutVec_63 : _GEN_4999; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_1_T_1 = 16'h3e + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_5002 = 6'h1 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5003 = 6'h2 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_2 : _GEN_5002; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5004 = 6'h3 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_3 : _GEN_5003; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5005 = 6'h4 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_4 : _GEN_5004; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5006 = 6'h5 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_5 : _GEN_5005; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5007 = 6'h6 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_6 : _GEN_5006; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5008 = 6'h7 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_7 : _GEN_5007; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5009 = 6'h8 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_8 : _GEN_5008; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5010 = 6'h9 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_9 : _GEN_5009; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5011 = 6'ha == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_10 : _GEN_5010; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5012 = 6'hb == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_11 : _GEN_5011; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5013 = 6'hc == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_12 : _GEN_5012; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5014 = 6'hd == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_13 : _GEN_5013; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5015 = 6'he == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_14 : _GEN_5014; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5016 = 6'hf == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_15 : _GEN_5015; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5017 = 6'h10 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_16 : _GEN_5016; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5018 = 6'h11 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_17 : _GEN_5017; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5019 = 6'h12 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_18 : _GEN_5018; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5020 = 6'h13 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_19 : _GEN_5019; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5021 = 6'h14 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_20 : _GEN_5020; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5022 = 6'h15 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_21 : _GEN_5021; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5023 = 6'h16 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_22 : _GEN_5022; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5024 = 6'h17 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_23 : _GEN_5023; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5025 = 6'h18 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_24 : _GEN_5024; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5026 = 6'h19 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_25 : _GEN_5025; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5027 = 6'h1a == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_26 : _GEN_5026; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5028 = 6'h1b == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_27 : _GEN_5027; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5029 = 6'h1c == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_28 : _GEN_5028; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5030 = 6'h1d == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_29 : _GEN_5029; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5031 = 6'h1e == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_30 : _GEN_5030; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5032 = 6'h1f == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_31 : _GEN_5031; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5033 = 6'h20 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_32 : _GEN_5032; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5034 = 6'h21 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_33 : _GEN_5033; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5035 = 6'h22 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_34 : _GEN_5034; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5036 = 6'h23 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_35 : _GEN_5035; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5037 = 6'h24 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_36 : _GEN_5036; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5038 = 6'h25 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_37 : _GEN_5037; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5039 = 6'h26 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_38 : _GEN_5038; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5040 = 6'h27 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_39 : _GEN_5039; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5041 = 6'h28 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_40 : _GEN_5040; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5042 = 6'h29 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_41 : _GEN_5041; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5043 = 6'h2a == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_42 : _GEN_5042; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5044 = 6'h2b == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_43 : _GEN_5043; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5045 = 6'h2c == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_44 : _GEN_5044; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5046 = 6'h2d == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_45 : _GEN_5045; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5047 = 6'h2e == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_46 : _GEN_5046; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5048 = 6'h2f == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_47 : _GEN_5047; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5049 = 6'h30 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_48 : _GEN_5048; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5050 = 6'h31 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_49 : _GEN_5049; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5051 = 6'h32 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_50 : _GEN_5050; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5052 = 6'h33 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_51 : _GEN_5051; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5053 = 6'h34 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_52 : _GEN_5052; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5054 = 6'h35 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_53 : _GEN_5053; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5055 = 6'h36 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_54 : _GEN_5054; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5056 = 6'h37 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_55 : _GEN_5055; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5057 = 6'h38 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_56 : _GEN_5056; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5058 = 6'h39 == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_57 : _GEN_5057; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5059 = 6'h3a == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_58 : _GEN_5058; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5060 = 6'h3b == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_59 : _GEN_5059; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5061 = 6'h3c == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_60 : _GEN_5060; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5062 = 6'h3d == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_61 : _GEN_5061; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5063 = 6'h3e == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_62 : _GEN_5062; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_1 = 6'h3f == _myHhdoutVec2_1_T_1[5:0] ? myHhdoutVec_63 : _GEN_5063; // @[hh_core.scala 149:{52,52}]
  wire [15:0] _myHhdoutVec2_0_T_1 = 16'h3f + io_hh_cnt; // @[hh_core.scala 149:72]
  wire [31:0] _GEN_5066 = 6'h1 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_1 : myHhdoutVec_0; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5067 = 6'h2 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_2 : _GEN_5066; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5068 = 6'h3 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_3 : _GEN_5067; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5069 = 6'h4 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_4 : _GEN_5068; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5070 = 6'h5 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_5 : _GEN_5069; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5071 = 6'h6 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_6 : _GEN_5070; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5072 = 6'h7 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_7 : _GEN_5071; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5073 = 6'h8 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_8 : _GEN_5072; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5074 = 6'h9 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_9 : _GEN_5073; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5075 = 6'ha == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_10 : _GEN_5074; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5076 = 6'hb == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_11 : _GEN_5075; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5077 = 6'hc == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_12 : _GEN_5076; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5078 = 6'hd == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_13 : _GEN_5077; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5079 = 6'he == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_14 : _GEN_5078; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5080 = 6'hf == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_15 : _GEN_5079; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5081 = 6'h10 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_16 : _GEN_5080; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5082 = 6'h11 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_17 : _GEN_5081; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5083 = 6'h12 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_18 : _GEN_5082; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5084 = 6'h13 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_19 : _GEN_5083; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5085 = 6'h14 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_20 : _GEN_5084; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5086 = 6'h15 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_21 : _GEN_5085; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5087 = 6'h16 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_22 : _GEN_5086; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5088 = 6'h17 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_23 : _GEN_5087; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5089 = 6'h18 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_24 : _GEN_5088; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5090 = 6'h19 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_25 : _GEN_5089; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5091 = 6'h1a == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_26 : _GEN_5090; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5092 = 6'h1b == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_27 : _GEN_5091; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5093 = 6'h1c == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_28 : _GEN_5092; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5094 = 6'h1d == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_29 : _GEN_5093; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5095 = 6'h1e == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_30 : _GEN_5094; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5096 = 6'h1f == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_31 : _GEN_5095; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5097 = 6'h20 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_32 : _GEN_5096; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5098 = 6'h21 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_33 : _GEN_5097; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5099 = 6'h22 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_34 : _GEN_5098; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5100 = 6'h23 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_35 : _GEN_5099; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5101 = 6'h24 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_36 : _GEN_5100; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5102 = 6'h25 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_37 : _GEN_5101; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5103 = 6'h26 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_38 : _GEN_5102; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5104 = 6'h27 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_39 : _GEN_5103; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5105 = 6'h28 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_40 : _GEN_5104; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5106 = 6'h29 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_41 : _GEN_5105; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5107 = 6'h2a == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_42 : _GEN_5106; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5108 = 6'h2b == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_43 : _GEN_5107; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5109 = 6'h2c == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_44 : _GEN_5108; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5110 = 6'h2d == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_45 : _GEN_5109; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5111 = 6'h2e == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_46 : _GEN_5110; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5112 = 6'h2f == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_47 : _GEN_5111; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5113 = 6'h30 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_48 : _GEN_5112; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5114 = 6'h31 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_49 : _GEN_5113; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5115 = 6'h32 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_50 : _GEN_5114; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5116 = 6'h33 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_51 : _GEN_5115; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5117 = 6'h34 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_52 : _GEN_5116; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5118 = 6'h35 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_53 : _GEN_5117; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5119 = 6'h36 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_54 : _GEN_5118; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5120 = 6'h37 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_55 : _GEN_5119; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5121 = 6'h38 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_56 : _GEN_5120; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5122 = 6'h39 == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_57 : _GEN_5121; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5123 = 6'h3a == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_58 : _GEN_5122; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5124 = 6'h3b == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_59 : _GEN_5123; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5125 = 6'h3c == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_60 : _GEN_5124; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5126 = 6'h3d == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_61 : _GEN_5125; // @[hh_core.scala 149:{52,52}]
  wire [31:0] _GEN_5127 = 6'h3e == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_62 : _GEN_5126; // @[hh_core.scala 149:{52,52}]
  wire [31:0] myHhdoutVec2_0 = 6'h3f == _myHhdoutVec2_0_T_1[5:0] ? myHhdoutVec_63 : _GEN_5127; // @[hh_core.scala 149:{52,52}]
  wire [255:0] myHhdoutWire_lo_lo_lo = {myHhdoutVec2_7,myHhdoutVec2_6,myHhdoutVec2_5,myHhdoutVec2_4,myHhdoutVec2_3,
    myHhdoutVec2_2,myHhdoutVec2_1,myHhdoutVec2_0}; // @[hh_core.scala 153:42]
  wire [511:0] myHhdoutWire_lo_lo = {myHhdoutVec2_15,myHhdoutVec2_14,myHhdoutVec2_13,myHhdoutVec2_12,myHhdoutVec2_11,
    myHhdoutVec2_10,myHhdoutVec2_9,myHhdoutVec2_8,myHhdoutWire_lo_lo_lo}; // @[hh_core.scala 153:42]
  wire [1023:0] myHhdoutWire_lo = {myHhdoutVec2_31,myHhdoutVec2_30,myHhdoutVec2_29,myHhdoutVec2_28,myHhdoutVec2_27,
    myHhdoutVec2_26,myHhdoutVec2_25,myHhdoutVec2_24,myHhdoutWire_lo_hi_lo,myHhdoutWire_lo_lo}; // @[hh_core.scala 153:42]
  wire [2047:0] myHhdoutWire = {myHhdoutWire_hi,myHhdoutWire_lo}; // @[hh_core.scala 153:42]
  wire [2047:0] _hh_dout_update_T_1 = myHhdoutWire >> _hh_din_update_T; // @[hh_core.scala 158:48]
  wire [2047:0] _GEN_5129 = io_hh_st ? _hh_dout_update_T_1 : hh_din_reg; // @[hh_core.scala 157:33 158:32 160:32]
  wire [2047:0] hh_dout = u_hh_datapath_io_hh_dout; // @[hh_core.scala 221:21 77:27]
  simple_dual simple_dual ( // @[hh_core.scala 163:31]
    .io_clka(simple_dual_io_clka),
    .io_clkb(simple_dual_io_clkb),
    .io_ena(simple_dual_io_ena),
    .io_enb(simple_dual_io_enb),
    .io_wea(simple_dual_io_wea),
    .io_addra(simple_dual_io_addra),
    .io_addrb(simple_dual_io_addrb),
    .io_dina(simple_dual_io_dina),
    .io_doutb(simple_dual_io_doutb)
  );
  simple_dual simple_dual_1 ( // @[hh_core.scala 175:31]
    .io_clka(simple_dual_1_io_clka),
    .io_clkb(simple_dual_1_io_clkb),
    .io_ena(simple_dual_1_io_ena),
    .io_enb(simple_dual_1_io_enb),
    .io_wea(simple_dual_1_io_wea),
    .io_addra(simple_dual_1_io_addra),
    .io_addrb(simple_dual_1_io_addrb),
    .io_dina(simple_dual_1_io_dina),
    .io_doutb(simple_dual_1_io_doutb)
  );
  simple_dual simple_dual_2 ( // @[hh_core.scala 186:31]
    .io_clka(simple_dual_2_io_clka),
    .io_clkb(simple_dual_2_io_clkb),
    .io_ena(simple_dual_2_io_ena),
    .io_enb(simple_dual_2_io_enb),
    .io_wea(simple_dual_2_io_wea),
    .io_addra(simple_dual_2_io_addra),
    .io_addrb(simple_dual_2_io_addrb),
    .io_dina(simple_dual_2_io_dina),
    .io_doutb(simple_dual_2_io_doutb)
  );
  hh_datapath_1 u_hh_datapath ( // @[hh_core.scala 197:38]
    .io_clk(u_hh_datapath_io_clk),
    .io_rst(u_hh_datapath_io_rst),
    .io_hh_cnt(u_hh_datapath_io_hh_cnt),
    .io_d1_rdy(u_hh_datapath_io_d1_rdy),
    .io_d1_vld(u_hh_datapath_io_d1_vld),
    .io_d2_vld(u_hh_datapath_io_d2_vld),
    .io_vk1_vld(u_hh_datapath_io_vk1_vld),
    .io_d3_rdy(u_hh_datapath_io_d3_rdy),
    .io_d3_vld(u_hh_datapath_io_d3_vld),
    .io_tk_vld(u_hh_datapath_io_tk_vld),
    .io_d4_rdy(u_hh_datapath_io_d4_rdy),
    .io_d5_rdy(u_hh_datapath_io_d5_rdy),
    .io_d5_vld(u_hh_datapath_io_d5_vld),
    .io_yj_sft(u_hh_datapath_io_yj_sft),
    .io_d4_sft(u_hh_datapath_io_d4_sft),
    .io_hh_din(u_hh_datapath_io_hh_din),
    .io_hh_dout(u_hh_datapath_io_hh_dout)
  );
  assign io_dmx0_mem_doutb = simple_dual_io_doutb; // @[hh_core.scala 173:31]
  assign io_dmx1_mem_doutb = simple_dual_1_io_doutb; // @[hh_core.scala 184:31]
  assign io_rtri_mem_doutb = simple_dual_2_io_doutb; // @[hh_core.scala 195:31]
  assign io_hh_dout = io_rst ? 2048'h0 : hh_dout; // @[hh_core.scala 222:25 223:27 225:24]
  assign simple_dual_io_clka = io_clk; // @[hh_core.scala 165:25]
  assign simple_dual_io_clkb = io_clk; // @[hh_core.scala 170:25]
  assign simple_dual_io_ena = io_dmx0_mem_ena; // @[hh_core.scala 166:24]
  assign simple_dual_io_enb = io_dmx0_mem_enb; // @[hh_core.scala 171:24]
  assign simple_dual_io_wea = io_dmx0_mem_wea; // @[hh_core.scala 167:24]
  assign simple_dual_io_addra = io_dmx0_mem_addra; // @[hh_core.scala 168:26]
  assign simple_dual_io_addrb = io_dmx0_mem_addrb; // @[hh_core.scala 172:26]
  assign simple_dual_io_dina = io_dmx0_mem_dina; // @[hh_core.scala 169:25]
  assign simple_dual_1_io_clka = io_clk; // @[hh_core.scala 176:25]
  assign simple_dual_1_io_clkb = io_clk; // @[hh_core.scala 181:25]
  assign simple_dual_1_io_ena = io_dmx1_mem_ena; // @[hh_core.scala 177:24]
  assign simple_dual_1_io_enb = io_dmx1_mem_enb; // @[hh_core.scala 182:24]
  assign simple_dual_1_io_wea = io_dmx1_mem_wea; // @[hh_core.scala 178:24]
  assign simple_dual_1_io_addra = io_dmx1_mem_addra; // @[hh_core.scala 179:26]
  assign simple_dual_1_io_addrb = io_dmx1_mem_addrb; // @[hh_core.scala 183:26]
  assign simple_dual_1_io_dina = io_dmx1_mem_dina; // @[hh_core.scala 180:25]
  assign simple_dual_2_io_clka = io_clk; // @[hh_core.scala 187:25]
  assign simple_dual_2_io_clkb = io_clk; // @[hh_core.scala 192:25]
  assign simple_dual_2_io_ena = io_rtri_mem_ena; // @[hh_core.scala 188:24]
  assign simple_dual_2_io_enb = io_rtri_mem_enb; // @[hh_core.scala 193:24]
  assign simple_dual_2_io_wea = io_rtri_mem_wea; // @[hh_core.scala 189:24]
  assign simple_dual_2_io_addra = io_rtri_mem_addra; // @[hh_core.scala 190:26]
  assign simple_dual_2_io_addrb = io_rtri_mem_addrb; // @[hh_core.scala 194:26]
  assign simple_dual_2_io_dina = io_rtri_mem_dina; // @[hh_core.scala 191:25]
  assign u_hh_datapath_io_clk = io_clk; // @[hh_core.scala 199:34]
  assign u_hh_datapath_io_rst = io_rst; // @[hh_core.scala 200:34]
  assign u_hh_datapath_io_hh_cnt = io_hh_cnt; // @[hh_core.scala 201:37]
  assign u_hh_datapath_io_d1_rdy = io_d1_rdy; // @[hh_core.scala 202:37]
  assign u_hh_datapath_io_d1_vld = io_d1_vld; // @[hh_core.scala 203:37]
  assign u_hh_datapath_io_d2_vld = io_d2_vld; // @[hh_core.scala 205:37]
  assign u_hh_datapath_io_vk1_vld = io_vk1_vld; // @[hh_core.scala 207:38]
  assign u_hh_datapath_io_d3_rdy = io_d3_rdy; // @[hh_core.scala 208:37]
  assign u_hh_datapath_io_d3_vld = io_d3_vld; // @[hh_core.scala 209:37]
  assign u_hh_datapath_io_tk_vld = io_tk_vld; // @[hh_core.scala 211:37]
  assign u_hh_datapath_io_d4_rdy = io_d4_rdy; // @[hh_core.scala 212:37]
  assign u_hh_datapath_io_d5_rdy = io_d5_rdy; // @[hh_core.scala 214:37]
  assign u_hh_datapath_io_d5_vld = io_d5_vld; // @[hh_core.scala 215:37]
  assign u_hh_datapath_io_yj_sft = io_yj_sft; // @[hh_core.scala 218:37]
  assign u_hh_datapath_io_d4_sft = io_d4_sft; // @[hh_core.scala 219:37]
  assign u_hh_datapath_io_hh_din = hh_din; // @[hh_core.scala 220:37]
  always @(posedge io_clk) begin
    if (io_rst) begin // @[hh_core.scala 87:25]
      hh0_din_rdy <= 1'h0; // @[hh_core.scala 88:29]
    end else begin
      hh0_din_rdy <= io_dmx0_mem_enb & io_rtri_mem_enb; // @[hh_core.scala 93:29]
    end
    if (io_rst) begin // @[hh_core.scala 87:25]
      hh1_din_rdy <= 1'h0; // @[hh_core.scala 89:29]
    end else begin
      hh1_din_rdy <= io_dmx1_mem_enb & io_rtri_mem_enb; // @[hh_core.scala 94:29]
    end
    if (io_rst) begin // @[hh_core.scala 87:25]
      hh_din_reg <= 2048'h0; // @[hh_core.scala 90:28]
    end else if (hh0_din_rdy | hh1_din_rdy) begin // @[hh_core.scala 100:44]
      if (_T) begin // @[hh_core.scala 133:44]
        hh_din_reg <= _hh_din_update_T_2; // @[hh_core.scala 134:31]
      end else if (io_rst) begin // @[hh_core.scala 135:31]
        hh_din_reg <= 2048'h0; // @[hh_core.scala 136:31]
      end
    end else if (io_hh_st) begin // @[hh_core.scala 102:33]
      if (io_rst) begin // @[hh_core.scala 155:25]
        hh_din_reg <= 2048'h0; // @[hh_core.scala 156:32]
      end else begin
        hh_din_reg <= _GEN_5129;
      end
    end
    if (io_rst) begin // @[hh_core.scala 87:25]
      hh_din <= 2048'h0; // @[hh_core.scala 90:28]
    end else if (hh0_din_rdy | hh1_din_rdy) begin // @[hh_core.scala 100:44]
      if (_T) begin // @[hh_core.scala 133:44]
        hh_din <= _hh_din_update_T_2; // @[hh_core.scala 134:31]
      end else if (io_rst) begin // @[hh_core.scala 135:31]
        hh_din <= 2048'h0; // @[hh_core.scala 136:31]
      end else begin
        hh_din <= hh_din_reg; // @[hh_core.scala 138:31]
      end
    end else if (io_hh_st) begin // @[hh_core.scala 102:33]
      if (io_rst) begin // @[hh_core.scala 155:25]
        hh_din <= 2048'h0; // @[hh_core.scala 156:32]
      end else begin
        hh_din <= _GEN_5129;
      end
    end else begin
      hh_din <= hh_din_reg; // @[hh_core.scala 106:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  hh0_din_rdy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hh1_din_rdy = _RAND_1[0:0];
  _RAND_2 = {64{`RANDOM}};
  hh_din_reg = _RAND_2[2047:0];
  _RAND_3 = {64{`RANDOM}};
  hh_din = _RAND_3[2047:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module tsqr_mc(
  input           clk,
  input           rst,
  input           tsqr_en,
  input  [15:0]   tile_no,
  input  [5:0]    dma_mem_ena,
  input  [127:0]  dma_mem_wea,
  input  [4:0]    dma_mem_addra,
  input  [1023:0] dma_mem_dina,
  input  [5:0]    dma_mem_enb,
  input  [4:0]    dma_mem_addrb,
  output [1023:0] dma_mem_doutb,
  output          mem0_fi_c_0,
  output          mem0_fi_c_1,
  output          mem1_fi_c_0,
  output          mem1_fi_c_1,
  output          tsqr_fi
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  fsms_0_clk; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_rst; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_tsqr_en; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_0_tile_no; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_0_hh_cnt; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_0_mx_cnt; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d1_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d1_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d2_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_vk1_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d3_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d3_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_tk_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d4_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d5_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d5_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_yj_sft; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_d4_sft; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_hh_st; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_mem0_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_mem1_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_tsqr_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_dmx0_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_0_dmx0_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_dmx0_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_dmx0_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_dmx0_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_dmx1_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_0_dmx1_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_dmx1_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_dmx1_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_dmx1_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_rtri_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_0_rtri_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_rtri_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_0_rtri_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_0_rtri_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_clk; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_rst; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_tsqr_en; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_1_tile_no; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_1_hh_cnt; // @[tsqr_mc.scala 1806:46]
  wire [15:0] fsms_1_mx_cnt; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d1_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d1_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d2_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_vk1_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d3_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d3_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_tk_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d4_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d5_rdy; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d5_vld; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_yj_sft; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_d4_sft; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_hh_st; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_mem0_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_mem1_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_tsqr_fi; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_dmx0_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_1_dmx0_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_dmx0_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_dmx0_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_dmx0_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_dmx1_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_1_dmx1_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_dmx1_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_dmx1_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_dmx1_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_rtri_mem_ena; // @[tsqr_mc.scala 1806:46]
  wire [127:0] fsms_1_rtri_mem_wea; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_rtri_mem_addra; // @[tsqr_mc.scala 1806:46]
  wire  fsms_1_rtri_mem_enb; // @[tsqr_mc.scala 1806:46]
  wire [4:0] fsms_1_rtri_mem_addrb; // @[tsqr_mc.scala 1806:46]
  wire  hh_core_io_clk; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_rst; // @[tsqr_mc.scala 1807:47]
  wire [15:0] hh_core_io_hh_cnt; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d1_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d1_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d2_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_vk1_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d3_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d3_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_tk_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d4_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d5_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d5_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_yj_sft; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_d4_sft; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_hh_st; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_dmx0_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_io_dmx0_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_dmx0_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_dmx0_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_dmx0_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_dmx0_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_dmx0_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_dmx1_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_io_dmx1_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_dmx1_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_dmx1_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_dmx1_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_dmx1_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_dmx1_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_rtri_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_io_rtri_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_rtri_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_rtri_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_io_rtri_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_io_rtri_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_io_rtri_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire [2047:0] hh_core_io_hh_dout; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_clk; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_rst; // @[tsqr_mc.scala 1807:47]
  wire [15:0] hh_core_1_io_hh_cnt; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d1_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d1_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d2_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_vk1_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d3_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d3_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_tk_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d4_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d5_rdy; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d5_vld; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_yj_sft; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_d4_sft; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_hh_st; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_dmx0_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_1_io_dmx0_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_dmx0_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_dmx0_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_dmx0_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_dmx0_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_dmx0_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_dmx1_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_1_io_dmx1_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_dmx1_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_dmx1_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_dmx1_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_dmx1_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_dmx1_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_rtri_mem_ena; // @[tsqr_mc.scala 1807:47]
  wire [127:0] hh_core_1_io_rtri_mem_wea; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_rtri_mem_addra; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_rtri_mem_dina; // @[tsqr_mc.scala 1807:47]
  wire  hh_core_1_io_rtri_mem_enb; // @[tsqr_mc.scala 1807:47]
  wire [4:0] hh_core_1_io_rtri_mem_addrb; // @[tsqr_mc.scala 1807:47]
  wire [1023:0] hh_core_1_io_rtri_mem_doutb; // @[tsqr_mc.scala 1807:47]
  wire [2047:0] hh_core_1_io_hh_dout; // @[tsqr_mc.scala 1807:47]
  reg  tsqr_fi_level_c_1; // @[tsqr_mc.scala 200:30]
  wire  _GEN_0 = tsqr_fi ? 1'h0 : tsqr_fi_level_c_1; // @[tsqr_mc.scala 207:28 200:30 208:32]
  wire  tsqr_fi_c_1 = fsms_1_tsqr_fi; // @[tsqr_mc.scala 175:26 1838:22]
  wire  _GEN_1 = tsqr_fi_c_1 | _GEN_0; // @[tsqr_mc.scala 205:33 206:32]
  wire  tsqr_en_c_1 = tsqr_en & ~tsqr_fi_level_c_1; // @[tsqr_mc.scala 215:34]
  wire [15:0] _tile_no_c_0_T = tile_no / 2'h2; // @[tsqr_mc.scala 224:48]
  wire [15:0] _tile_no_c_0_T_2 = _tile_no_c_0_T - 16'h1; // @[tsqr_mc.scala 224:62]
  wire [15:0] _tile_no_c_0_T_4 = _tile_no_c_0_T_2 + 16'h1; // @[tsqr_mc.scala 224:67]
  wire  tsqr_fi_c_0 = fsms_0_tsqr_fi; // @[tsqr_mc.scala 175:26 1838:22]
  wire  fsm_rtri_mem_ena_c_0 = fsms_0_rtri_mem_ena; // @[tsqr_mc.scala 1849:31 186:35]
  wire  fsm_rtri_mem_ena_c_1 = fsms_1_rtri_mem_ena; // @[tsqr_mc.scala 1849:31 186:35]
  wire  rtri_mem_ena_c_1 = dma_mem_ena[2] | fsm_rtri_mem_ena_c_1; // @[tsqr_mc.scala 252:68]
  wire  fsm_dmx0_mem_ena_c_0 = fsms_0_dmx0_mem_ena; // @[tsqr_mc.scala 176:35 1839:31]
  wire [15:0] mx_cnt_c_1 = fsms_1_mx_cnt; // @[tsqr_mc.scala 154:25 1816:21]
  wire [15:0] _wr_dmx0_mem_ena_0_T_2 = _tile_no_c_0_T - 16'h2; // @[tsqr_mc.scala 1783:97]
  wire  _wr_dmx0_mem_ena_0_T_4 = rtri_mem_ena_c_1 & mx_cnt_c_1 == _wr_dmx0_mem_ena_0_T_2; // @[tsqr_mc.scala 1783:56]
  wire  wr_dmx0_mem_ena_0 = rtri_mem_ena_c_1 & mx_cnt_c_1 == _wr_dmx0_mem_ena_0_T_2 & tile_no[1]; // @[tsqr_mc.scala 1783:103]
  wire  fsm_dmx0_mem_ena_c_1 = fsms_1_dmx0_mem_ena; // @[tsqr_mc.scala 176:35 1839:31]
  wire  fsm_dmx1_mem_ena_c_0 = fsms_0_dmx1_mem_ena; // @[tsqr_mc.scala 181:35 1844:31]
  wire  wr_dmx1_mem_ena_0 = _wr_dmx0_mem_ena_0_T_4 & ~tile_no[1]; // @[tsqr_mc.scala 1782:103]
  wire  fsm_dmx1_mem_ena_c_1 = fsms_1_dmx1_mem_ena; // @[tsqr_mc.scala 181:35 1844:31]
  wire [127:0] fsm_rtri_mem_wea_c_0 = fsms_0_rtri_mem_wea; // @[tsqr_mc.scala 1850:31 187:35]
  wire [127:0] fsm_rtri_mem_wea_c_1 = fsms_1_rtri_mem_wea; // @[tsqr_mc.scala 1850:31 187:35]
  wire [127:0] _GEN_8 = wr_dmx0_mem_ena_0 ? fsm_rtri_mem_wea_c_1 : 128'h0; // @[tsqr_mc.scala 372:53 373:45 375:45]
  wire [127:0] fsm_dmx0_mem_wea_c_0 = fsms_0_dmx0_mem_wea; // @[tsqr_mc.scala 177:35 1840:31]
  wire [127:0] _GEN_9 = fsm_dmx0_mem_ena_c_0 ? fsm_dmx0_mem_wea_c_0 : _GEN_8; // @[tsqr_mc.scala 370:56 371:45]
  wire [127:0] fsm_dmx0_mem_wea_c_1 = fsms_1_dmx0_mem_wea; // @[tsqr_mc.scala 177:35 1840:31]
  wire [127:0] _GEN_12 = wr_dmx1_mem_ena_0 ? fsm_rtri_mem_wea_c_1 : 128'h0; // @[tsqr_mc.scala 594:53 595:45 597:45]
  wire [127:0] fsm_dmx1_mem_wea_c_0 = fsms_0_dmx1_mem_wea; // @[tsqr_mc.scala 182:35 1845:31]
  wire [127:0] _GEN_13 = fsm_dmx1_mem_ena_c_0 ? fsm_dmx1_mem_wea_c_0 : _GEN_12; // @[tsqr_mc.scala 592:56 593:45]
  wire [127:0] fsm_dmx1_mem_wea_c_1 = fsms_1_dmx1_mem_wea; // @[tsqr_mc.scala 182:35 1845:31]
  wire [4:0] fsm_rtri_mem_addra_c_0 = fsms_0_rtri_mem_addra; // @[tsqr_mc.scala 1851:33 188:37]
  wire [4:0] fsm_rtri_mem_addra_c_1 = fsms_1_rtri_mem_addra; // @[tsqr_mc.scala 1851:33 188:37]
  wire [4:0] _GEN_18 = wr_dmx0_mem_ena_0 ? fsm_rtri_mem_addra_c_1 : 5'h0; // @[tsqr_mc.scala 830:53 831:47 833:47]
  wire [4:0] fsm_dmx0_mem_addra_c_0 = fsms_0_dmx0_mem_addra; // @[tsqr_mc.scala 178:37 1841:33]
  wire [4:0] _GEN_19 = fsm_dmx0_mem_ena_c_0 ? fsm_dmx0_mem_addra_c_0 : _GEN_18; // @[tsqr_mc.scala 828:56 829:47]
  wire [4:0] fsm_dmx0_mem_addra_c_1 = fsms_1_dmx0_mem_addra; // @[tsqr_mc.scala 178:37 1841:33]
  wire [4:0] _GEN_22 = wr_dmx1_mem_ena_0 ? fsm_rtri_mem_addra_c_1 : 5'h0; // @[tsqr_mc.scala 1052:53 1053:47 1055:47]
  wire [4:0] fsm_dmx1_mem_addra_c_0 = fsms_0_dmx1_mem_addra; // @[tsqr_mc.scala 183:37 1846:33]
  wire [4:0] _GEN_23 = fsm_dmx1_mem_ena_c_0 ? fsm_dmx1_mem_addra_c_0 : _GEN_22; // @[tsqr_mc.scala 1050:56 1051:47]
  wire [4:0] fsm_dmx1_mem_addra_c_1 = fsms_1_dmx1_mem_addra; // @[tsqr_mc.scala 183:37 1846:33]
  wire [2047:0] hh_dout_c_0 = hh_core_io_hh_dout; // @[tsqr_mc.scala 1897:22 191:26]
  wire [1023:0] _GEN_26 = fsm_rtri_mem_ena_c_0 ? hh_dout_c_0[2047:1024] : 1024'h0; // @[tsqr_mc.scala 1261:42 1262:32 1264:32]
  wire [2047:0] hh_dout_c_1 = hh_core_1_io_hh_dout; // @[tsqr_mc.scala 1897:22 191:26]
  wire [1023:0] _GEN_28 = fsm_rtri_mem_ena_c_1 ? hh_dout_c_1[2047:1024] : 1024'h0; // @[tsqr_mc.scala 1261:42 1262:32 1264:32]
  wire [1023:0] _GEN_30 = wr_dmx0_mem_ena_0 ? hh_dout_c_1[2047:1024] : 1024'h0; // @[tsqr_mc.scala 1294:53 1295:46 1297:46]
  wire [1023:0] _GEN_31 = fsm_dmx0_mem_ena_c_0 ? hh_dout_c_0[1023:0] : _GEN_30; // @[tsqr_mc.scala 1292:56 1293:46]
  wire [1023:0] _GEN_33 = fsm_dmx0_mem_ena_c_1 ? hh_dout_c_1[1023:0] : 1024'h0; // @[tsqr_mc.scala 1274:48 1275:38 1277:38]
  wire [1023:0] _GEN_35 = wr_dmx1_mem_ena_0 ? hh_dout_c_1[2047:1024] : 1024'h0; // @[tsqr_mc.scala 1520:53 1521:46 1523:46]
  wire [1023:0] _GEN_36 = fsm_dmx1_mem_ena_c_0 ? hh_dout_c_0[1023:0] : _GEN_35; // @[tsqr_mc.scala 1518:56 1519:46]
  wire [1023:0] _GEN_38 = fsm_dmx1_mem_ena_c_1 ? hh_dout_c_1[1023:0] : 1024'h0; // @[tsqr_mc.scala 1500:48 1501:38 1503:38]
  wire  fsm_rtri_mem_enb_c_0 = fsms_0_rtri_mem_enb; // @[tsqr_mc.scala 1852:31 189:35]
  wire  fsm_dmx0_mem_enb_c_0 = fsms_0_dmx0_mem_enb; // @[tsqr_mc.scala 179:35 1842:31]
  wire  fsm_dmx1_mem_enb_c_0 = fsms_0_dmx1_mem_enb; // @[tsqr_mc.scala 184:35 1847:31]
  wire  fsm_rtri_mem_enb_c_1 = fsms_1_rtri_mem_enb; // @[tsqr_mc.scala 1852:31 189:35]
  wire  fsm_dmx0_mem_enb_c_1 = fsms_1_dmx0_mem_enb; // @[tsqr_mc.scala 179:35 1842:31]
  wire  fsm_dmx1_mem_enb_c_1 = fsms_1_dmx1_mem_enb; // @[tsqr_mc.scala 184:35 1847:31]
  wire [4:0] fsm_rtri_mem_addrb_c_0 = fsms_0_rtri_mem_addrb; // @[tsqr_mc.scala 1853:33 190:37]
  wire [4:0] fsm_rtri_mem_addrb_c_1 = fsms_1_rtri_mem_addrb; // @[tsqr_mc.scala 1853:33 190:37]
  wire [4:0] fsm_dmx0_mem_addrb_c_0 = fsms_0_dmx0_mem_addrb; // @[tsqr_mc.scala 180:37 1843:33]
  wire [4:0] fsm_dmx0_mem_addrb_c_1 = fsms_1_dmx0_mem_addrb; // @[tsqr_mc.scala 180:37 1843:33]
  wire [4:0] fsm_dmx1_mem_addrb_c_0 = fsms_0_dmx1_mem_addrb; // @[tsqr_mc.scala 1848:33 185:37]
  wire [4:0] fsm_dmx1_mem_addrb_c_1 = fsms_1_dmx1_mem_addrb; // @[tsqr_mc.scala 1848:33 185:37]
  wire [5:0] _T_30 = dma_mem_enb[5] ? 6'h20 : 6'h0; // @[Mux.scala 47:70]
  wire [5:0] _T_31 = dma_mem_enb[4] ? 6'h10 : _T_30; // @[Mux.scala 47:70]
  wire [5:0] _T_32 = dma_mem_enb[3] ? 6'h8 : _T_31; // @[Mux.scala 47:70]
  wire [5:0] _T_33 = dma_mem_enb[2] ? 6'h4 : _T_32; // @[Mux.scala 47:70]
  wire [5:0] _T_34 = dma_mem_enb[1] ? 6'h2 : _T_33; // @[Mux.scala 47:70]
  wire [5:0] _T_35 = dma_mem_enb[0] ? 6'h1 : _T_34; // @[Mux.scala 47:70]
  wire [5:0] _dma_mem_doutb_T_13 = _T_35 + 6'h3; // @[tsqr_mc.scala 1775:93]
  wire [5:0] _dma_mem_doutb_T_14 = _dma_mem_doutb_T_13 / 2'h3; // @[tsqr_mc.scala 1775:99]
  wire [5:0] _dma_mem_doutb_T_16 = 6'h2 - _dma_mem_doutb_T_14; // @[tsqr_mc.scala 1775:59]
  wire [1023:0] dmx1_mem_doutb_c_0 = hh_core_io_dmx1_mem_doutb; // @[tsqr_mc.scala 1765:32 1900:29]
  wire [1023:0] dmx1_mem_doutb_c_1 = hh_core_1_io_dmx1_mem_doutb; // @[tsqr_mc.scala 1765:32 1900:29]
  wire [1023:0] _GEN_47 = _dma_mem_doutb_T_16[0] ? dmx1_mem_doutb_c_1 : dmx1_mem_doutb_c_0; // @[tsqr_mc.scala 1775:{27,27}]
  fsm fsms_0 ( // @[tsqr_mc.scala 1806:46]
    .clk(fsms_0_clk),
    .rst(fsms_0_rst),
    .tsqr_en(fsms_0_tsqr_en),
    .tile_no(fsms_0_tile_no),
    .hh_cnt(fsms_0_hh_cnt),
    .mx_cnt(fsms_0_mx_cnt),
    .d1_rdy(fsms_0_d1_rdy),
    .d1_vld(fsms_0_d1_vld),
    .d2_vld(fsms_0_d2_vld),
    .vk1_vld(fsms_0_vk1_vld),
    .d3_rdy(fsms_0_d3_rdy),
    .d3_vld(fsms_0_d3_vld),
    .tk_vld(fsms_0_tk_vld),
    .d4_rdy(fsms_0_d4_rdy),
    .d5_rdy(fsms_0_d5_rdy),
    .d5_vld(fsms_0_d5_vld),
    .yj_sft(fsms_0_yj_sft),
    .d4_sft(fsms_0_d4_sft),
    .hh_st(fsms_0_hh_st),
    .mem0_fi(fsms_0_mem0_fi),
    .mem1_fi(fsms_0_mem1_fi),
    .tsqr_fi(fsms_0_tsqr_fi),
    .dmx0_mem_ena(fsms_0_dmx0_mem_ena),
    .dmx0_mem_wea(fsms_0_dmx0_mem_wea),
    .dmx0_mem_addra(fsms_0_dmx0_mem_addra),
    .dmx0_mem_enb(fsms_0_dmx0_mem_enb),
    .dmx0_mem_addrb(fsms_0_dmx0_mem_addrb),
    .dmx1_mem_ena(fsms_0_dmx1_mem_ena),
    .dmx1_mem_wea(fsms_0_dmx1_mem_wea),
    .dmx1_mem_addra(fsms_0_dmx1_mem_addra),
    .dmx1_mem_enb(fsms_0_dmx1_mem_enb),
    .dmx1_mem_addrb(fsms_0_dmx1_mem_addrb),
    .rtri_mem_ena(fsms_0_rtri_mem_ena),
    .rtri_mem_wea(fsms_0_rtri_mem_wea),
    .rtri_mem_addra(fsms_0_rtri_mem_addra),
    .rtri_mem_enb(fsms_0_rtri_mem_enb),
    .rtri_mem_addrb(fsms_0_rtri_mem_addrb)
  );
  fsm fsms_1 ( // @[tsqr_mc.scala 1806:46]
    .clk(fsms_1_clk),
    .rst(fsms_1_rst),
    .tsqr_en(fsms_1_tsqr_en),
    .tile_no(fsms_1_tile_no),
    .hh_cnt(fsms_1_hh_cnt),
    .mx_cnt(fsms_1_mx_cnt),
    .d1_rdy(fsms_1_d1_rdy),
    .d1_vld(fsms_1_d1_vld),
    .d2_vld(fsms_1_d2_vld),
    .vk1_vld(fsms_1_vk1_vld),
    .d3_rdy(fsms_1_d3_rdy),
    .d3_vld(fsms_1_d3_vld),
    .tk_vld(fsms_1_tk_vld),
    .d4_rdy(fsms_1_d4_rdy),
    .d5_rdy(fsms_1_d5_rdy),
    .d5_vld(fsms_1_d5_vld),
    .yj_sft(fsms_1_yj_sft),
    .d4_sft(fsms_1_d4_sft),
    .hh_st(fsms_1_hh_st),
    .mem0_fi(fsms_1_mem0_fi),
    .mem1_fi(fsms_1_mem1_fi),
    .tsqr_fi(fsms_1_tsqr_fi),
    .dmx0_mem_ena(fsms_1_dmx0_mem_ena),
    .dmx0_mem_wea(fsms_1_dmx0_mem_wea),
    .dmx0_mem_addra(fsms_1_dmx0_mem_addra),
    .dmx0_mem_enb(fsms_1_dmx0_mem_enb),
    .dmx0_mem_addrb(fsms_1_dmx0_mem_addrb),
    .dmx1_mem_ena(fsms_1_dmx1_mem_ena),
    .dmx1_mem_wea(fsms_1_dmx1_mem_wea),
    .dmx1_mem_addra(fsms_1_dmx1_mem_addra),
    .dmx1_mem_enb(fsms_1_dmx1_mem_enb),
    .dmx1_mem_addrb(fsms_1_dmx1_mem_addrb),
    .rtri_mem_ena(fsms_1_rtri_mem_ena),
    .rtri_mem_wea(fsms_1_rtri_mem_wea),
    .rtri_mem_addra(fsms_1_rtri_mem_addra),
    .rtri_mem_enb(fsms_1_rtri_mem_enb),
    .rtri_mem_addrb(fsms_1_rtri_mem_addrb)
  );
  hh_core hh_core ( // @[tsqr_mc.scala 1807:47]
    .io_clk(hh_core_io_clk),
    .io_rst(hh_core_io_rst),
    .io_hh_cnt(hh_core_io_hh_cnt),
    .io_d1_rdy(hh_core_io_d1_rdy),
    .io_d1_vld(hh_core_io_d1_vld),
    .io_d2_vld(hh_core_io_d2_vld),
    .io_vk1_vld(hh_core_io_vk1_vld),
    .io_d3_rdy(hh_core_io_d3_rdy),
    .io_d3_vld(hh_core_io_d3_vld),
    .io_tk_vld(hh_core_io_tk_vld),
    .io_d4_rdy(hh_core_io_d4_rdy),
    .io_d5_rdy(hh_core_io_d5_rdy),
    .io_d5_vld(hh_core_io_d5_vld),
    .io_yj_sft(hh_core_io_yj_sft),
    .io_d4_sft(hh_core_io_d4_sft),
    .io_hh_st(hh_core_io_hh_st),
    .io_dmx0_mem_ena(hh_core_io_dmx0_mem_ena),
    .io_dmx0_mem_wea(hh_core_io_dmx0_mem_wea),
    .io_dmx0_mem_addra(hh_core_io_dmx0_mem_addra),
    .io_dmx0_mem_dina(hh_core_io_dmx0_mem_dina),
    .io_dmx0_mem_enb(hh_core_io_dmx0_mem_enb),
    .io_dmx0_mem_addrb(hh_core_io_dmx0_mem_addrb),
    .io_dmx0_mem_doutb(hh_core_io_dmx0_mem_doutb),
    .io_dmx1_mem_ena(hh_core_io_dmx1_mem_ena),
    .io_dmx1_mem_wea(hh_core_io_dmx1_mem_wea),
    .io_dmx1_mem_addra(hh_core_io_dmx1_mem_addra),
    .io_dmx1_mem_dina(hh_core_io_dmx1_mem_dina),
    .io_dmx1_mem_enb(hh_core_io_dmx1_mem_enb),
    .io_dmx1_mem_addrb(hh_core_io_dmx1_mem_addrb),
    .io_dmx1_mem_doutb(hh_core_io_dmx1_mem_doutb),
    .io_rtri_mem_ena(hh_core_io_rtri_mem_ena),
    .io_rtri_mem_wea(hh_core_io_rtri_mem_wea),
    .io_rtri_mem_addra(hh_core_io_rtri_mem_addra),
    .io_rtri_mem_dina(hh_core_io_rtri_mem_dina),
    .io_rtri_mem_enb(hh_core_io_rtri_mem_enb),
    .io_rtri_mem_addrb(hh_core_io_rtri_mem_addrb),
    .io_rtri_mem_doutb(hh_core_io_rtri_mem_doutb),
    .io_hh_dout(hh_core_io_hh_dout)
  );
  hh_core hh_core_1 ( // @[tsqr_mc.scala 1807:47]
    .io_clk(hh_core_1_io_clk),
    .io_rst(hh_core_1_io_rst),
    .io_hh_cnt(hh_core_1_io_hh_cnt),
    .io_d1_rdy(hh_core_1_io_d1_rdy),
    .io_d1_vld(hh_core_1_io_d1_vld),
    .io_d2_vld(hh_core_1_io_d2_vld),
    .io_vk1_vld(hh_core_1_io_vk1_vld),
    .io_d3_rdy(hh_core_1_io_d3_rdy),
    .io_d3_vld(hh_core_1_io_d3_vld),
    .io_tk_vld(hh_core_1_io_tk_vld),
    .io_d4_rdy(hh_core_1_io_d4_rdy),
    .io_d5_rdy(hh_core_1_io_d5_rdy),
    .io_d5_vld(hh_core_1_io_d5_vld),
    .io_yj_sft(hh_core_1_io_yj_sft),
    .io_d4_sft(hh_core_1_io_d4_sft),
    .io_hh_st(hh_core_1_io_hh_st),
    .io_dmx0_mem_ena(hh_core_1_io_dmx0_mem_ena),
    .io_dmx0_mem_wea(hh_core_1_io_dmx0_mem_wea),
    .io_dmx0_mem_addra(hh_core_1_io_dmx0_mem_addra),
    .io_dmx0_mem_dina(hh_core_1_io_dmx0_mem_dina),
    .io_dmx0_mem_enb(hh_core_1_io_dmx0_mem_enb),
    .io_dmx0_mem_addrb(hh_core_1_io_dmx0_mem_addrb),
    .io_dmx0_mem_doutb(hh_core_1_io_dmx0_mem_doutb),
    .io_dmx1_mem_ena(hh_core_1_io_dmx1_mem_ena),
    .io_dmx1_mem_wea(hh_core_1_io_dmx1_mem_wea),
    .io_dmx1_mem_addra(hh_core_1_io_dmx1_mem_addra),
    .io_dmx1_mem_dina(hh_core_1_io_dmx1_mem_dina),
    .io_dmx1_mem_enb(hh_core_1_io_dmx1_mem_enb),
    .io_dmx1_mem_addrb(hh_core_1_io_dmx1_mem_addrb),
    .io_dmx1_mem_doutb(hh_core_1_io_dmx1_mem_doutb),
    .io_rtri_mem_ena(hh_core_1_io_rtri_mem_ena),
    .io_rtri_mem_wea(hh_core_1_io_rtri_mem_wea),
    .io_rtri_mem_addra(hh_core_1_io_rtri_mem_addra),
    .io_rtri_mem_dina(hh_core_1_io_rtri_mem_dina),
    .io_rtri_mem_enb(hh_core_1_io_rtri_mem_enb),
    .io_rtri_mem_addrb(hh_core_1_io_rtri_mem_addrb),
    .io_rtri_mem_doutb(hh_core_1_io_rtri_mem_doutb),
    .io_hh_dout(hh_core_1_io_hh_dout)
  );
  assign dma_mem_doutb = rst ? 1024'h0 : _GEN_47; // @[tsqr_mc.scala 1767:14 1768:23 1775:27]
  assign mem0_fi_c_0 = fsms_0_mem0_fi; // @[tsqr_mc.scala 1836:22]
  assign mem0_fi_c_1 = fsms_1_mem0_fi; // @[tsqr_mc.scala 1836:22]
  assign mem1_fi_c_0 = fsms_0_mem1_fi; // @[tsqr_mc.scala 1837:22]
  assign mem1_fi_c_1 = fsms_1_mem1_fi; // @[tsqr_mc.scala 1837:22]
  assign tsqr_fi = tsqr_en & tsqr_fi_c_0; // @[tsqr_mc.scala 244:23 245:17 247:17]
  assign fsms_0_clk = clk; // @[tsqr_mc.scala 1811:21]
  assign fsms_0_rst = rst; // @[tsqr_mc.scala 1812:21]
  assign fsms_0_tsqr_en = tsqr_en; // @[tsqr_mc.scala 215:34]
  assign fsms_0_tile_no = tsqr_en ? _tile_no_c_0_T_4 : 16'h0; // @[tsqr_mc.scala 219:29 224:36 240:28]
  assign fsms_1_clk = clk; // @[tsqr_mc.scala 1811:21]
  assign fsms_1_rst = rst; // @[tsqr_mc.scala 1812:21]
  assign fsms_1_tsqr_en = tsqr_en & ~tsqr_fi_level_c_1; // @[tsqr_mc.scala 215:34]
  assign fsms_1_tile_no = tsqr_en_c_1 ? _tile_no_c_0_T_2 : 16'h0; // @[tsqr_mc.scala 219:29 221:32 240:28]
  assign hh_core_io_clk = clk; // @[tsqr_mc.scala 1855:22]
  assign hh_core_io_rst = rst; // @[tsqr_mc.scala 1856:22]
  assign hh_core_io_hh_cnt = fsms_0_hh_cnt; // @[tsqr_mc.scala 155:25 1815:21]
  assign hh_core_io_d1_rdy = fsms_0_d1_rdy; // @[tsqr_mc.scala 156:25 1817:21]
  assign hh_core_io_d1_vld = fsms_0_d1_vld; // @[tsqr_mc.scala 157:25 1818:21]
  assign hh_core_io_d2_vld = fsms_0_d2_vld; // @[tsqr_mc.scala 159:25 1820:21]
  assign hh_core_io_vk1_vld = fsms_0_vk1_vld; // @[tsqr_mc.scala 161:26 1822:22]
  assign hh_core_io_d3_rdy = fsms_0_d3_rdy; // @[tsqr_mc.scala 162:25 1823:21]
  assign hh_core_io_d3_vld = fsms_0_d3_vld; // @[tsqr_mc.scala 163:25 1824:21]
  assign hh_core_io_tk_vld = fsms_0_tk_vld; // @[tsqr_mc.scala 165:25 1826:21]
  assign hh_core_io_d4_rdy = fsms_0_d4_rdy; // @[tsqr_mc.scala 166:25 1827:21]
  assign hh_core_io_d5_rdy = fsms_0_d5_rdy; // @[tsqr_mc.scala 168:25 1829:21]
  assign hh_core_io_d5_vld = fsms_0_d5_vld; // @[tsqr_mc.scala 169:25 1830:21]
  assign hh_core_io_yj_sft = fsms_0_yj_sft; // @[tsqr_mc.scala 172:25 1833:21]
  assign hh_core_io_d4_sft = fsms_0_d4_sft; // @[tsqr_mc.scala 173:25 1834:21]
  assign hh_core_io_hh_st = fsms_0_hh_st; // @[tsqr_mc.scala 174:24 1835:20]
  assign hh_core_io_dmx0_mem_ena = dma_mem_ena[4] | fsm_dmx0_mem_ena_c_0 | wr_dmx0_mem_ena_0; // @[tsqr_mc.scala 265:114]
  assign hh_core_io_dmx0_mem_wea = dma_mem_ena[4] ? dma_mem_wea : _GEN_9; // @[tsqr_mc.scala 368:61 369:45]
  assign hh_core_io_dmx0_mem_addra = dma_mem_ena[4] ? dma_mem_addra : _GEN_19; // @[tsqr_mc.scala 826:61 827:47]
  assign hh_core_io_dmx0_mem_dina = dma_mem_ena[4] ? dma_mem_dina : _GEN_31; // @[tsqr_mc.scala 1290:61 1291:46]
  assign hh_core_io_dmx0_mem_enb = dma_mem_enb[4] | fsm_dmx0_mem_enb_c_0; // @[tsqr_mc.scala 1728:68]
  assign hh_core_io_dmx0_mem_addrb = dma_mem_ena[4] ? dma_mem_addrb : fsm_dmx0_mem_addrb_c_0; // @[tsqr_mc.scala 1747:50 1748:33 1750:33]
  assign hh_core_io_dmx1_mem_ena = dma_mem_ena[3] | fsm_dmx1_mem_ena_c_0 | wr_dmx1_mem_ena_0; // @[tsqr_mc.scala 307:106]
  assign hh_core_io_dmx1_mem_wea = dma_mem_ena[3] ? dma_mem_wea : _GEN_13; // @[tsqr_mc.scala 590:59 591:45]
  assign hh_core_io_dmx1_mem_addra = dma_mem_ena[3] ? dma_mem_addra : _GEN_23; // @[tsqr_mc.scala 1048:59 1049:47]
  assign hh_core_io_dmx1_mem_dina = dma_mem_ena[3] ? dma_mem_dina : _GEN_36; // @[tsqr_mc.scala 1516:59 1517:46]
  assign hh_core_io_dmx1_mem_enb = dma_mem_enb[3] | fsm_dmx1_mem_enb_c_0; // @[tsqr_mc.scala 1729:70]
  assign hh_core_io_dmx1_mem_addrb = dma_mem_ena[3] ? dma_mem_addrb : fsm_dmx1_mem_addrb_c_0; // @[tsqr_mc.scala 1755:52 1756:33 1758:33]
  assign hh_core_io_rtri_mem_ena = dma_mem_ena[5] | fsm_rtri_mem_ena_c_0; // @[tsqr_mc.scala 252:68]
  assign hh_core_io_rtri_mem_wea = dma_mem_ena[5] ? dma_mem_wea : fsm_rtri_mem_wea_c_0; // @[tsqr_mc.scala 343:50 344:31 346:31]
  assign hh_core_io_rtri_mem_addra = dma_mem_ena[5] ? dma_mem_addra : fsm_rtri_mem_addra_c_0; // @[tsqr_mc.scala 801:50 802:33 804:33]
  assign hh_core_io_rtri_mem_dina = dma_mem_ena[5] ? dma_mem_dina : _GEN_26; // @[tsqr_mc.scala 1259:50 1260:32]
  assign hh_core_io_rtri_mem_enb = dma_mem_enb[5] | fsm_rtri_mem_enb_c_0; // @[tsqr_mc.scala 1727:68]
  assign hh_core_io_rtri_mem_addrb = dma_mem_ena[5] ? dma_mem_addrb : fsm_rtri_mem_addrb_c_0; // @[tsqr_mc.scala 1739:50 1740:33 1742:33]
  assign hh_core_1_io_clk = clk; // @[tsqr_mc.scala 1855:22]
  assign hh_core_1_io_rst = rst; // @[tsqr_mc.scala 1856:22]
  assign hh_core_1_io_hh_cnt = fsms_1_hh_cnt; // @[tsqr_mc.scala 155:25 1815:21]
  assign hh_core_1_io_d1_rdy = fsms_1_d1_rdy; // @[tsqr_mc.scala 156:25 1817:21]
  assign hh_core_1_io_d1_vld = fsms_1_d1_vld; // @[tsqr_mc.scala 157:25 1818:21]
  assign hh_core_1_io_d2_vld = fsms_1_d2_vld; // @[tsqr_mc.scala 159:25 1820:21]
  assign hh_core_1_io_vk1_vld = fsms_1_vk1_vld; // @[tsqr_mc.scala 161:26 1822:22]
  assign hh_core_1_io_d3_rdy = fsms_1_d3_rdy; // @[tsqr_mc.scala 162:25 1823:21]
  assign hh_core_1_io_d3_vld = fsms_1_d3_vld; // @[tsqr_mc.scala 163:25 1824:21]
  assign hh_core_1_io_tk_vld = fsms_1_tk_vld; // @[tsqr_mc.scala 165:25 1826:21]
  assign hh_core_1_io_d4_rdy = fsms_1_d4_rdy; // @[tsqr_mc.scala 166:25 1827:21]
  assign hh_core_1_io_d5_rdy = fsms_1_d5_rdy; // @[tsqr_mc.scala 168:25 1829:21]
  assign hh_core_1_io_d5_vld = fsms_1_d5_vld; // @[tsqr_mc.scala 169:25 1830:21]
  assign hh_core_1_io_yj_sft = fsms_1_yj_sft; // @[tsqr_mc.scala 172:25 1833:21]
  assign hh_core_1_io_d4_sft = fsms_1_d4_sft; // @[tsqr_mc.scala 173:25 1834:21]
  assign hh_core_1_io_hh_st = fsms_1_hh_st; // @[tsqr_mc.scala 174:24 1835:20]
  assign hh_core_1_io_dmx0_mem_ena = dma_mem_ena[1] | fsm_dmx0_mem_ena_c_1; // @[tsqr_mc.scala 259:80]
  assign hh_core_1_io_dmx0_mem_wea = dma_mem_ena[1] ? dma_mem_wea : fsm_dmx0_mem_wea_c_1; // @[tsqr_mc.scala 354:54 355:37 357:37]
  assign hh_core_1_io_dmx0_mem_addra = dma_mem_ena[1] ? dma_mem_addra : fsm_dmx0_mem_addra_c_1; // @[tsqr_mc.scala 812:54 813:39 815:39]
  assign hh_core_1_io_dmx0_mem_dina = dma_mem_ena[1] ? dma_mem_dina : _GEN_33; // @[tsqr_mc.scala 1272:56 1273:38]
  assign hh_core_1_io_dmx0_mem_enb = dma_mem_enb[1] | fsm_dmx0_mem_enb_c_1; // @[tsqr_mc.scala 1728:68]
  assign hh_core_1_io_dmx0_mem_addrb = dma_mem_ena[1] ? dma_mem_addrb : fsm_dmx0_mem_addrb_c_1; // @[tsqr_mc.scala 1747:50 1748:33 1750:33]
  assign hh_core_1_io_dmx1_mem_ena = dma_mem_ena[0] | fsm_dmx1_mem_ena_c_1; // @[tsqr_mc.scala 301:72]
  assign hh_core_1_io_dmx1_mem_wea = dma_mem_ena[0] ? dma_mem_wea : fsm_dmx1_mem_wea_c_1; // @[tsqr_mc.scala 576:52 577:37 579:37]
  assign hh_core_1_io_dmx1_mem_addra = dma_mem_ena[0] ? dma_mem_addra : fsm_dmx1_mem_addra_c_1; // @[tsqr_mc.scala 1034:52 1035:39 1037:39]
  assign hh_core_1_io_dmx1_mem_dina = dma_mem_ena[0] ? dma_mem_dina : _GEN_38; // @[tsqr_mc.scala 1498:52 1499:38]
  assign hh_core_1_io_dmx1_mem_enb = dma_mem_enb[0] | fsm_dmx1_mem_enb_c_1; // @[tsqr_mc.scala 1729:70]
  assign hh_core_1_io_dmx1_mem_addrb = dma_mem_ena[0] ? dma_mem_addrb : fsm_dmx1_mem_addrb_c_1; // @[tsqr_mc.scala 1755:52 1756:33 1758:33]
  assign hh_core_1_io_rtri_mem_ena = dma_mem_ena[2] | fsm_rtri_mem_ena_c_1; // @[tsqr_mc.scala 252:68]
  assign hh_core_1_io_rtri_mem_wea = dma_mem_ena[2] ? dma_mem_wea : fsm_rtri_mem_wea_c_1; // @[tsqr_mc.scala 343:50 344:31 346:31]
  assign hh_core_1_io_rtri_mem_addra = dma_mem_ena[2] ? dma_mem_addra : fsm_rtri_mem_addra_c_1; // @[tsqr_mc.scala 801:50 802:33 804:33]
  assign hh_core_1_io_rtri_mem_dina = dma_mem_ena[2] ? dma_mem_dina : _GEN_28; // @[tsqr_mc.scala 1259:50 1260:32]
  assign hh_core_1_io_rtri_mem_enb = dma_mem_enb[2] | fsm_rtri_mem_enb_c_1; // @[tsqr_mc.scala 1727:68]
  assign hh_core_1_io_rtri_mem_addrb = dma_mem_ena[2] ? dma_mem_addrb : fsm_rtri_mem_addrb_c_1; // @[tsqr_mc.scala 1739:50 1740:33 1742:33]
  always @(posedge clk) begin
    if (rst) begin // @[tsqr_mc.scala 203:18]
      tsqr_fi_level_c_1 <= 1'h0; // @[tsqr_mc.scala 204:32]
    end else begin
      tsqr_fi_level_c_1 <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tsqr_fi_level_c_1 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

