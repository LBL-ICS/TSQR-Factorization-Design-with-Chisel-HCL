`ifdef ST_WIDTH_INF_16
reg [31:0] golden_yjp0  ;
reg [31:0] golden_yjp1  ;
reg [31:0] golden_yjp2  ;
reg [31:0] golden_yjp3  ;
reg [31:0] golden_yjp4  ;
reg [31:0] golden_yjp5  ;
reg [31:0] golden_yjp6  ;
reg [31:0] golden_yjp7  ;
reg [31:0] golden_yjp8  ;
reg [31:0] golden_yjp9  ;
reg [31:0] golden_yjp10 ;
reg [31:0] golden_yjp11 ;
reg [31:0] golden_yjp12 ;
reg [31:0] golden_yjp13 ;
reg [31:0] golden_yjp14 ;
reg [31:0] golden_yjp15 ;
`endif //ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32 
reg [31:0] golden_yjp16 ;
reg [31:0] golden_yjp17 ;
reg [31:0] golden_yjp18 ;
reg [31:0] golden_yjp19 ;
reg [31:0] golden_yjp20 ;
reg [31:0] golden_yjp21 ;
reg [31:0] golden_yjp22 ;
reg [31:0] golden_yjp23 ;
reg [31:0] golden_yjp24 ;
reg [31:0] golden_yjp25 ;
reg [31:0] golden_yjp26 ;
reg [31:0] golden_yjp27 ;
reg [31:0] golden_yjp28 ;
reg [31:0] golden_yjp29 ;
reg [31:0] golden_yjp30 ;
reg [31:0] golden_yjp31 ;
`endif //ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64 
reg [31:0] golden_yjp32 ;
reg [31:0] golden_yjp33 ;
reg [31:0] golden_yjp34 ;
reg [31:0] golden_yjp35 ;
reg [31:0] golden_yjp36 ;
reg [31:0] golden_yjp37 ;
reg [31:0] golden_yjp38 ;
reg [31:0] golden_yjp39 ;
reg [31:0] golden_yjp40 ;
reg [31:0] golden_yjp41 ;
reg [31:0] golden_yjp42 ;
reg [31:0] golden_yjp43 ;
reg [31:0] golden_yjp44 ;
reg [31:0] golden_yjp45 ;
reg [31:0] golden_yjp46 ;
reg [31:0] golden_yjp47 ;
reg [31:0] golden_yjp48 ;
reg [31:0] golden_yjp49 ;
reg [31:0] golden_yjp50 ;
reg [31:0] golden_yjp51 ;
reg [31:0] golden_yjp52 ;
reg [31:0] golden_yjp53 ;
reg [31:0] golden_yjp54 ;
reg [31:0] golden_yjp55 ;
reg [31:0] golden_yjp56 ;
reg [31:0] golden_yjp57 ;
reg [31:0] golden_yjp58 ;
reg [31:0] golden_yjp59 ;
reg [31:0] golden_yjp60 ;
reg [31:0] golden_yjp61 ;
reg [31:0] golden_yjp62 ;
reg [31:0] golden_yjp63 ;
`endif //ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128 
reg [31:0] golden_yjp64 ;
reg [31:0] golden_yjp65 ;
reg [31:0] golden_yjp66 ;
reg [31:0] golden_yjp67 ;
reg [31:0] golden_yjp68 ;
reg [31:0] golden_yjp69 ;
reg [31:0] golden_yjp70 ;
reg [31:0] golden_yjp71 ;
reg [31:0] golden_yjp72 ;
reg [31:0] golden_yjp73 ;
reg [31:0] golden_yjp74 ;
reg [31:0] golden_yjp75 ;
reg [31:0] golden_yjp76 ;
reg [31:0] golden_yjp77 ;
reg [31:0] golden_yjp78 ;
reg [31:0] golden_yjp79 ;
reg [31:0] golden_yjp80 ;
reg [31:0] golden_yjp81 ;
reg [31:0] golden_yjp82 ;
reg [31:0] golden_yjp83 ;
reg [31:0] golden_yjp84 ;
reg [31:0] golden_yjp85 ;
reg [31:0] golden_yjp86 ;
reg [31:0] golden_yjp87 ;
reg [31:0] golden_yjp88 ;
reg [31:0] golden_yjp89 ;
reg [31:0] golden_yjp90 ;
reg [31:0] golden_yjp91 ;
reg [31:0] golden_yjp92 ;
reg [31:0] golden_yjp93 ;
reg [31:0] golden_yjp94 ;
reg [31:0] golden_yjp95 ;
reg [31:0] golden_yjp96 ;
reg [31:0] golden_yjp97 ;
reg [31:0] golden_yjp98 ;
reg [31:0] golden_yjp99 ;
reg [31:0] golden_yjp100;
reg [31:0] golden_yjp101;
reg [31:0] golden_yjp102;
reg [31:0] golden_yjp103;
reg [31:0] golden_yjp104;
reg [31:0] golden_yjp105;
reg [31:0] golden_yjp106;
reg [31:0] golden_yjp107;
reg [31:0] golden_yjp108;
reg [31:0] golden_yjp109;
reg [31:0] golden_yjp110;
reg [31:0] golden_yjp111;
reg [31:0] golden_yjp112;
reg [31:0] golden_yjp113;
reg [31:0] golden_yjp114;
reg [31:0] golden_yjp115;
reg [31:0] golden_yjp116;
reg [31:0] golden_yjp117;
reg [31:0] golden_yjp118;
reg [31:0] golden_yjp119;
reg [31:0] golden_yjp120;
reg [31:0] golden_yjp121;
reg [31:0] golden_yjp122;
reg [31:0] golden_yjp123;
reg [31:0] golden_yjp124;
reg [31:0] golden_yjp125;
reg [31:0] golden_yjp126;
reg [31:0] golden_yjp127;
`endif //ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256 
reg [31:0] golden_yjp128;
reg [31:0] golden_yjp129;
reg [31:0] golden_yjp130;
reg [31:0] golden_yjp131;
reg [31:0] golden_yjp132;
reg [31:0] golden_yjp133;
reg [31:0] golden_yjp134;
reg [31:0] golden_yjp135;
reg [31:0] golden_yjp136;
reg [31:0] golden_yjp137;
reg [31:0] golden_yjp138;
reg [31:0] golden_yjp139;
reg [31:0] golden_yjp140;
reg [31:0] golden_yjp141;
reg [31:0] golden_yjp142;
reg [31:0] golden_yjp143;
reg [31:0] golden_yjp144;
reg [31:0] golden_yjp145;
reg [31:0] golden_yjp146;
reg [31:0] golden_yjp147;
reg [31:0] golden_yjp148;
reg [31:0] golden_yjp149;
reg [31:0] golden_yjp150;
reg [31:0] golden_yjp151;
reg [31:0] golden_yjp152;
reg [31:0] golden_yjp153;
reg [31:0] golden_yjp154;
reg [31:0] golden_yjp155;
reg [31:0] golden_yjp156;
reg [31:0] golden_yjp157;
reg [31:0] golden_yjp158;
reg [31:0] golden_yjp159;
reg [31:0] golden_yjp160;
reg [31:0] golden_yjp161;
reg [31:0] golden_yjp162;
reg [31:0] golden_yjp163;
reg [31:0] golden_yjp164;
reg [31:0] golden_yjp165;
reg [31:0] golden_yjp166;
reg [31:0] golden_yjp167;
reg [31:0] golden_yjp168;
reg [31:0] golden_yjp169;
reg [31:0] golden_yjp170;
reg [31:0] golden_yjp171;
reg [31:0] golden_yjp172;
reg [31:0] golden_yjp173;
reg [31:0] golden_yjp174;
reg [31:0] golden_yjp175;
reg [31:0] golden_yjp176;
reg [31:0] golden_yjp177;
reg [31:0] golden_yjp178;
reg [31:0] golden_yjp179;
reg [31:0] golden_yjp180;
reg [31:0] golden_yjp181;
reg [31:0] golden_yjp182;
reg [31:0] golden_yjp183;
reg [31:0] golden_yjp184;
reg [31:0] golden_yjp185;
reg [31:0] golden_yjp186;
reg [31:0] golden_yjp187;
reg [31:0] golden_yjp188;
reg [31:0] golden_yjp189;
reg [31:0] golden_yjp190;
reg [31:0] golden_yjp191;
reg [31:0] golden_yjp192;
reg [31:0] golden_yjp193;
reg [31:0] golden_yjp194;
reg [31:0] golden_yjp195;
reg [31:0] golden_yjp196;
reg [31:0] golden_yjp197;
reg [31:0] golden_yjp198;
reg [31:0] golden_yjp199;
reg [31:0] golden_yjp200;
reg [31:0] golden_yjp201;
reg [31:0] golden_yjp202;
reg [31:0] golden_yjp203;
reg [31:0] golden_yjp204;
reg [31:0] golden_yjp205;
reg [31:0] golden_yjp206;
reg [31:0] golden_yjp207;
reg [31:0] golden_yjp208;
reg [31:0] golden_yjp209;
reg [31:0] golden_yjp210;
reg [31:0] golden_yjp211;
reg [31:0] golden_yjp212;
reg [31:0] golden_yjp213;
reg [31:0] golden_yjp214;
reg [31:0] golden_yjp215;
reg [31:0] golden_yjp216;
reg [31:0] golden_yjp217;
reg [31:0] golden_yjp218;
reg [31:0] golden_yjp219;
reg [31:0] golden_yjp220;
reg [31:0] golden_yjp221;
reg [31:0] golden_yjp222;
reg [31:0] golden_yjp223;
reg [31:0] golden_yjp224;
reg [31:0] golden_yjp225;
reg [31:0] golden_yjp226;
reg [31:0] golden_yjp227;
reg [31:0] golden_yjp228;
reg [31:0] golden_yjp229;
reg [31:0] golden_yjp230;
reg [31:0] golden_yjp231;
reg [31:0] golden_yjp232;
reg [31:0] golden_yjp233;
reg [31:0] golden_yjp234;
reg [31:0] golden_yjp235;
reg [31:0] golden_yjp236;
reg [31:0] golden_yjp237;
reg [31:0] golden_yjp238;
reg [31:0] golden_yjp239;
reg [31:0] golden_yjp240;
reg [31:0] golden_yjp241;
reg [31:0] golden_yjp242;
reg [31:0] golden_yjp243;
reg [31:0] golden_yjp244;
reg [31:0] golden_yjp245;
reg [31:0] golden_yjp246;
reg [31:0] golden_yjp247;
reg [31:0] golden_yjp248;
reg [31:0] golden_yjp249;
reg [31:0] golden_yjp250;
reg [31:0] golden_yjp251;
reg [31:0] golden_yjp252;
reg [31:0] golden_yjp253;
reg [31:0] golden_yjp254;
reg [31:0] golden_yjp255;
`endif //ST_WIDTH_INF_256
`ifdef ST_WIDTH_INF_16
reg [31:0] dut_yjp0     ;
reg [31:0] dut_yjp1     ;
reg [31:0] dut_yjp2     ;
reg [31:0] dut_yjp3     ;
reg [31:0] dut_yjp4     ;
reg [31:0] dut_yjp5     ;
reg [31:0] dut_yjp6     ;
reg [31:0] dut_yjp7     ;
reg [31:0] dut_yjp8     ;
reg [31:0] dut_yjp9     ;
reg [31:0] dut_yjp10    ;
reg [31:0] dut_yjp11    ;
reg [31:0] dut_yjp12    ;
reg [31:0] dut_yjp13    ;
reg [31:0] dut_yjp14    ;
reg [31:0] dut_yjp15    ;
`endif //ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32
reg [31:0] dut_yjp16    ;
reg [31:0] dut_yjp17    ;
reg [31:0] dut_yjp18    ;
reg [31:0] dut_yjp19    ;
reg [31:0] dut_yjp20    ;
reg [31:0] dut_yjp21    ;
reg [31:0] dut_yjp22    ;
reg [31:0] dut_yjp23    ;
reg [31:0] dut_yjp24    ;
reg [31:0] dut_yjp25    ;
reg [31:0] dut_yjp26    ;
reg [31:0] dut_yjp27    ;
reg [31:0] dut_yjp28    ;
reg [31:0] dut_yjp29    ;
reg [31:0] dut_yjp30    ;
reg [31:0] dut_yjp31    ;
`endif //ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64
reg [31:0] dut_yjp32    ;
reg [31:0] dut_yjp33    ;
reg [31:0] dut_yjp34    ;
reg [31:0] dut_yjp35    ;
reg [31:0] dut_yjp36    ;
reg [31:0] dut_yjp37    ;
reg [31:0] dut_yjp38    ;
reg [31:0] dut_yjp39    ;
reg [31:0] dut_yjp40    ;
reg [31:0] dut_yjp41    ;
reg [31:0] dut_yjp42    ;
reg [31:0] dut_yjp43    ;
reg [31:0] dut_yjp44    ;
reg [31:0] dut_yjp45    ;
reg [31:0] dut_yjp46    ;
reg [31:0] dut_yjp47    ;
reg [31:0] dut_yjp48    ;
reg [31:0] dut_yjp49    ;
reg [31:0] dut_yjp50    ;
reg [31:0] dut_yjp51    ;
reg [31:0] dut_yjp52    ;
reg [31:0] dut_yjp53    ;
reg [31:0] dut_yjp54    ;
reg [31:0] dut_yjp55    ;
reg [31:0] dut_yjp56    ;
reg [31:0] dut_yjp57    ;
reg [31:0] dut_yjp58    ;
reg [31:0] dut_yjp59    ;
reg [31:0] dut_yjp60    ;
reg [31:0] dut_yjp61    ;
reg [31:0] dut_yjp62    ;
reg [31:0] dut_yjp63    ;
`endif //ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128
reg [31:0] dut_yjp64    ;
reg [31:0] dut_yjp65    ;
reg [31:0] dut_yjp66    ;
reg [31:0] dut_yjp67    ;
reg [31:0] dut_yjp68    ;
reg [31:0] dut_yjp69    ;
reg [31:0] dut_yjp70    ;
reg [31:0] dut_yjp71    ;
reg [31:0] dut_yjp72    ;
reg [31:0] dut_yjp73    ;
reg [31:0] dut_yjp74    ;
reg [31:0] dut_yjp75    ;
reg [31:0] dut_yjp76    ;
reg [31:0] dut_yjp77    ;
reg [31:0] dut_yjp78    ;
reg [31:0] dut_yjp79    ;
reg [31:0] dut_yjp80    ;
reg [31:0] dut_yjp81    ;
reg [31:0] dut_yjp82    ;
reg [31:0] dut_yjp83    ;
reg [31:0] dut_yjp84    ;
reg [31:0] dut_yjp85    ;
reg [31:0] dut_yjp86    ;
reg [31:0] dut_yjp87    ;
reg [31:0] dut_yjp88    ;
reg [31:0] dut_yjp89    ;
reg [31:0] dut_yjp90    ;
reg [31:0] dut_yjp91    ;
reg [31:0] dut_yjp92    ;
reg [31:0] dut_yjp93    ;
reg [31:0] dut_yjp94    ;
reg [31:0] dut_yjp95    ;
reg [31:0] dut_yjp96    ;
reg [31:0] dut_yjp97    ;
reg [31:0] dut_yjp98    ;
reg [31:0] dut_yjp99    ;
reg [31:0] dut_yjp100   ;
reg [31:0] dut_yjp101   ;
reg [31:0] dut_yjp102   ;
reg [31:0] dut_yjp103   ;
reg [31:0] dut_yjp104   ;
reg [31:0] dut_yjp105   ;
reg [31:0] dut_yjp106   ;
reg [31:0] dut_yjp107   ;
reg [31:0] dut_yjp108   ;
reg [31:0] dut_yjp109   ;
reg [31:0] dut_yjp110   ;
reg [31:0] dut_yjp111   ;
reg [31:0] dut_yjp112   ;
reg [31:0] dut_yjp113   ;
reg [31:0] dut_yjp114   ;
reg [31:0] dut_yjp115   ;
reg [31:0] dut_yjp116   ;
reg [31:0] dut_yjp117   ;
reg [31:0] dut_yjp118   ;
reg [31:0] dut_yjp119   ;
reg [31:0] dut_yjp120   ;
reg [31:0] dut_yjp121   ;
reg [31:0] dut_yjp122   ;
reg [31:0] dut_yjp123   ;
reg [31:0] dut_yjp124   ;
reg [31:0] dut_yjp125   ;
reg [31:0] dut_yjp126   ;
reg [31:0] dut_yjp127   ;
`endif //ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256
reg [31:0] dut_yjp128   ;
reg [31:0] dut_yjp129   ;
reg [31:0] dut_yjp130   ;
reg [31:0] dut_yjp131   ;
reg [31:0] dut_yjp132   ;
reg [31:0] dut_yjp133   ;
reg [31:0] dut_yjp134   ;
reg [31:0] dut_yjp135   ;
reg [31:0] dut_yjp136   ;
reg [31:0] dut_yjp137   ;
reg [31:0] dut_yjp138   ;
reg [31:0] dut_yjp139   ;
reg [31:0] dut_yjp140   ;
reg [31:0] dut_yjp141   ;
reg [31:0] dut_yjp142   ;
reg [31:0] dut_yjp143   ;
reg [31:0] dut_yjp144   ;
reg [31:0] dut_yjp145   ;
reg [31:0] dut_yjp146   ;
reg [31:0] dut_yjp147   ;
reg [31:0] dut_yjp148   ;
reg [31:0] dut_yjp149   ;
reg [31:0] dut_yjp150   ;
reg [31:0] dut_yjp151   ;
reg [31:0] dut_yjp152   ;
reg [31:0] dut_yjp153   ;
reg [31:0] dut_yjp154   ;
reg [31:0] dut_yjp155   ;
reg [31:0] dut_yjp156   ;
reg [31:0] dut_yjp157   ;
reg [31:0] dut_yjp158   ;
reg [31:0] dut_yjp159   ;
reg [31:0] dut_yjp160   ;
reg [31:0] dut_yjp161   ;
reg [31:0] dut_yjp162   ;
reg [31:0] dut_yjp163   ;
reg [31:0] dut_yjp164   ;
reg [31:0] dut_yjp165   ;
reg [31:0] dut_yjp166   ;
reg [31:0] dut_yjp167   ;
reg [31:0] dut_yjp168   ;
reg [31:0] dut_yjp169   ;
reg [31:0] dut_yjp170   ;
reg [31:0] dut_yjp171   ;
reg [31:0] dut_yjp172   ;
reg [31:0] dut_yjp173   ;
reg [31:0] dut_yjp174   ;
reg [31:0] dut_yjp175   ;
reg [31:0] dut_yjp176   ;
reg [31:0] dut_yjp177   ;
reg [31:0] dut_yjp178   ;
reg [31:0] dut_yjp179   ;
reg [31:0] dut_yjp180   ;
reg [31:0] dut_yjp181   ;
reg [31:0] dut_yjp182   ;
reg [31:0] dut_yjp183   ;
reg [31:0] dut_yjp184   ;
reg [31:0] dut_yjp185   ;
reg [31:0] dut_yjp186   ;
reg [31:0] dut_yjp187   ;
reg [31:0] dut_yjp188   ;
reg [31:0] dut_yjp189   ;
reg [31:0] dut_yjp190   ;
reg [31:0] dut_yjp191   ;
reg [31:0] dut_yjp192   ;
reg [31:0] dut_yjp193   ;
reg [31:0] dut_yjp194   ;
reg [31:0] dut_yjp195   ;
reg [31:0] dut_yjp196   ;
reg [31:0] dut_yjp197   ;
reg [31:0] dut_yjp198   ;
reg [31:0] dut_yjp199   ;
reg [31:0] dut_yjp200   ;
reg [31:0] dut_yjp201   ;
reg [31:0] dut_yjp202   ;
reg [31:0] dut_yjp203   ;
reg [31:0] dut_yjp204   ;
reg [31:0] dut_yjp205   ;
reg [31:0] dut_yjp206   ;
reg [31:0] dut_yjp207   ;
reg [31:0] dut_yjp208   ;
reg [31:0] dut_yjp209   ;
reg [31:0] dut_yjp210   ;
reg [31:0] dut_yjp211   ;
reg [31:0] dut_yjp212   ;
reg [31:0] dut_yjp213   ;
reg [31:0] dut_yjp214   ;
reg [31:0] dut_yjp215   ;
reg [31:0] dut_yjp216   ;
reg [31:0] dut_yjp217   ;
reg [31:0] dut_yjp218   ;
reg [31:0] dut_yjp219   ;
reg [31:0] dut_yjp220   ;
reg [31:0] dut_yjp221   ;
reg [31:0] dut_yjp222   ;
reg [31:0] dut_yjp223   ;
reg [31:0] dut_yjp224   ;
reg [31:0] dut_yjp225   ;
reg [31:0] dut_yjp226   ;
reg [31:0] dut_yjp227   ;
reg [31:0] dut_yjp228   ;
reg [31:0] dut_yjp229   ;
reg [31:0] dut_yjp230   ;
reg [31:0] dut_yjp231   ;
reg [31:0] dut_yjp232   ;
reg [31:0] dut_yjp233   ;
reg [31:0] dut_yjp234   ;
reg [31:0] dut_yjp235   ;
reg [31:0] dut_yjp236   ;
reg [31:0] dut_yjp237   ;
reg [31:0] dut_yjp238   ;
reg [31:0] dut_yjp239   ;
reg [31:0] dut_yjp240   ;
reg [31:0] dut_yjp241   ;
reg [31:0] dut_yjp242   ;
reg [31:0] dut_yjp243   ;
reg [31:0] dut_yjp244   ;
reg [31:0] dut_yjp245   ;
reg [31:0] dut_yjp246   ;
reg [31:0] dut_yjp247   ;
reg [31:0] dut_yjp248   ;
reg [31:0] dut_yjp249   ;
reg [31:0] dut_yjp250   ;
reg [31:0] dut_yjp251   ;
reg [31:0] dut_yjp252   ;
reg [31:0] dut_yjp253   ;
reg [31:0] dut_yjp254   ;
reg [31:0] dut_yjp255   ;
`endif //ST_WIDTH_INF_256
`ifdef ST_WIDTH_INF_16
real golden_real_yjp0  ;
real golden_real_yjp1  ;
real golden_real_yjp2  ;
real golden_real_yjp3  ;
real golden_real_yjp4  ;
real golden_real_yjp5  ;
real golden_real_yjp6  ;
real golden_real_yjp7  ;
real golden_real_yjp8  ;
real golden_real_yjp9  ;
real golden_real_yjp10 ;
real golden_real_yjp11 ;
real golden_real_yjp12 ;
real golden_real_yjp13 ;
real golden_real_yjp14 ;
real golden_real_yjp15 ;
`endif //ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32 
real golden_real_yjp16 ;
real golden_real_yjp17 ;
real golden_real_yjp18 ;
real golden_real_yjp19 ;
real golden_real_yjp20 ;
real golden_real_yjp21 ;
real golden_real_yjp22 ;
real golden_real_yjp23 ;
real golden_real_yjp24 ;
real golden_real_yjp25 ;
real golden_real_yjp26 ;
real golden_real_yjp27 ;
real golden_real_yjp28 ;
real golden_real_yjp29 ;
real golden_real_yjp30 ;
real golden_real_yjp31 ;
`endif //ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64 
real golden_real_yjp32 ;
real golden_real_yjp33 ;
real golden_real_yjp34 ;
real golden_real_yjp35 ;
real golden_real_yjp36 ;
real golden_real_yjp37 ;
real golden_real_yjp38 ;
real golden_real_yjp39 ;
real golden_real_yjp40 ;
real golden_real_yjp41 ;
real golden_real_yjp42 ;
real golden_real_yjp43 ;
real golden_real_yjp44 ;
real golden_real_yjp45 ;
real golden_real_yjp46 ;
real golden_real_yjp47 ;
real golden_real_yjp48 ;
real golden_real_yjp49 ;
real golden_real_yjp50 ;
real golden_real_yjp51 ;
real golden_real_yjp52 ;
real golden_real_yjp53 ;
real golden_real_yjp54 ;
real golden_real_yjp55 ;
real golden_real_yjp56 ;
real golden_real_yjp57 ;
real golden_real_yjp58 ;
real golden_real_yjp59 ;
real golden_real_yjp60 ;
real golden_real_yjp61 ;
real golden_real_yjp62 ;
real golden_real_yjp63 ;
`endif //ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128 
real golden_real_yjp64 ;
real golden_real_yjp65 ;
real golden_real_yjp66 ;
real golden_real_yjp67 ;
real golden_real_yjp68 ;
real golden_real_yjp69 ;
real golden_real_yjp70 ;
real golden_real_yjp71 ;
real golden_real_yjp72 ;
real golden_real_yjp73 ;
real golden_real_yjp74 ;
real golden_real_yjp75 ;
real golden_real_yjp76 ;
real golden_real_yjp77 ;
real golden_real_yjp78 ;
real golden_real_yjp79 ;
real golden_real_yjp80 ;
real golden_real_yjp81 ;
real golden_real_yjp82 ;
real golden_real_yjp83 ;
real golden_real_yjp84 ;
real golden_real_yjp85 ;
real golden_real_yjp86 ;
real golden_real_yjp87 ;
real golden_real_yjp88 ;
real golden_real_yjp89 ;
real golden_real_yjp90 ;
real golden_real_yjp91 ;
real golden_real_yjp92 ;
real golden_real_yjp93 ;
real golden_real_yjp94 ;
real golden_real_yjp95 ;
real golden_real_yjp96 ;
real golden_real_yjp97 ;
real golden_real_yjp98 ;
real golden_real_yjp99 ;
real golden_real_yjp100;
real golden_real_yjp101;
real golden_real_yjp102;
real golden_real_yjp103;
real golden_real_yjp104;
real golden_real_yjp105;
real golden_real_yjp106;
real golden_real_yjp107;
real golden_real_yjp108;
real golden_real_yjp109;
real golden_real_yjp110;
real golden_real_yjp111;
real golden_real_yjp112;
real golden_real_yjp113;
real golden_real_yjp114;
real golden_real_yjp115;
real golden_real_yjp116;
real golden_real_yjp117;
real golden_real_yjp118;
real golden_real_yjp119;
real golden_real_yjp120;
real golden_real_yjp121;
real golden_real_yjp122;
real golden_real_yjp123;
real golden_real_yjp124;
real golden_real_yjp125;
real golden_real_yjp126;
real golden_real_yjp127;
`endif //ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256 
real golden_real_yjp128;
real golden_real_yjp129;
real golden_real_yjp130;
real golden_real_yjp131;
real golden_real_yjp132;
real golden_real_yjp133;
real golden_real_yjp134;
real golden_real_yjp135;
real golden_real_yjp136;
real golden_real_yjp137;
real golden_real_yjp138;
real golden_real_yjp139;
real golden_real_yjp140;
real golden_real_yjp141;
real golden_real_yjp142;
real golden_real_yjp143;
real golden_real_yjp144;
real golden_real_yjp145;
real golden_real_yjp146;
real golden_real_yjp147;
real golden_real_yjp148;
real golden_real_yjp149;
real golden_real_yjp150;
real golden_real_yjp151;
real golden_real_yjp152;
real golden_real_yjp153;
real golden_real_yjp154;
real golden_real_yjp155;
real golden_real_yjp156;
real golden_real_yjp157;
real golden_real_yjp158;
real golden_real_yjp159;
real golden_real_yjp160;
real golden_real_yjp161;
real golden_real_yjp162;
real golden_real_yjp163;
real golden_real_yjp164;
real golden_real_yjp165;
real golden_real_yjp166;
real golden_real_yjp167;
real golden_real_yjp168;
real golden_real_yjp169;
real golden_real_yjp170;
real golden_real_yjp171;
real golden_real_yjp172;
real golden_real_yjp173;
real golden_real_yjp174;
real golden_real_yjp175;
real golden_real_yjp176;
real golden_real_yjp177;
real golden_real_yjp178;
real golden_real_yjp179;
real golden_real_yjp180;
real golden_real_yjp181;
real golden_real_yjp182;
real golden_real_yjp183;
real golden_real_yjp184;
real golden_real_yjp185;
real golden_real_yjp186;
real golden_real_yjp187;
real golden_real_yjp188;
real golden_real_yjp189;
real golden_real_yjp190;
real golden_real_yjp191;
real golden_real_yjp192;
real golden_real_yjp193;
real golden_real_yjp194;
real golden_real_yjp195;
real golden_real_yjp196;
real golden_real_yjp197;
real golden_real_yjp198;
real golden_real_yjp199;
real golden_real_yjp200;
real golden_real_yjp201;
real golden_real_yjp202;
real golden_real_yjp203;
real golden_real_yjp204;
real golden_real_yjp205;
real golden_real_yjp206;
real golden_real_yjp207;
real golden_real_yjp208;
real golden_real_yjp209;
real golden_real_yjp210;
real golden_real_yjp211;
real golden_real_yjp212;
real golden_real_yjp213;
real golden_real_yjp214;
real golden_real_yjp215;
real golden_real_yjp216;
real golden_real_yjp217;
real golden_real_yjp218;
real golden_real_yjp219;
real golden_real_yjp220;
real golden_real_yjp221;
real golden_real_yjp222;
real golden_real_yjp223;
real golden_real_yjp224;
real golden_real_yjp225;
real golden_real_yjp226;
real golden_real_yjp227;
real golden_real_yjp228;
real golden_real_yjp229;
real golden_real_yjp230;
real golden_real_yjp231;
real golden_real_yjp232;
real golden_real_yjp233;
real golden_real_yjp234;
real golden_real_yjp235;
real golden_real_yjp236;
real golden_real_yjp237;
real golden_real_yjp238;
real golden_real_yjp239;
real golden_real_yjp240;
real golden_real_yjp241;
real golden_real_yjp242;
real golden_real_yjp243;
real golden_real_yjp244;
real golden_real_yjp245;
real golden_real_yjp246;
real golden_real_yjp247;
real golden_real_yjp248;
real golden_real_yjp249;
real golden_real_yjp250;
real golden_real_yjp251;
real golden_real_yjp252;
real golden_real_yjp253;
real golden_real_yjp254;
real golden_real_yjp255;
`endif //ST_WIDTH_INF_256
`ifdef ST_WIDTH_INF_16
real dut_real_yjp0     ;
real dut_real_yjp1     ;
real dut_real_yjp2     ;
real dut_real_yjp3     ;
real dut_real_yjp4     ;
real dut_real_yjp5     ;
real dut_real_yjp6     ;
real dut_real_yjp7     ;
real dut_real_yjp8     ;
real dut_real_yjp9     ;
real dut_real_yjp10    ;
real dut_real_yjp11    ;
real dut_real_yjp12    ;
real dut_real_yjp13    ;
real dut_real_yjp14    ;
real dut_real_yjp15    ;
`endif //ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32
real dut_real_yjp16    ;
real dut_real_yjp17    ;
real dut_real_yjp18    ;
real dut_real_yjp19    ;
real dut_real_yjp20    ;
real dut_real_yjp21    ;
real dut_real_yjp22    ;
real dut_real_yjp23    ;
real dut_real_yjp24    ;
real dut_real_yjp25    ;
real dut_real_yjp26    ;
real dut_real_yjp27    ;
real dut_real_yjp28    ;
real dut_real_yjp29    ;
real dut_real_yjp30    ;
real dut_real_yjp31    ;
`endif //ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64
real dut_real_yjp32    ;
real dut_real_yjp33    ;
real dut_real_yjp34    ;
real dut_real_yjp35    ;
real dut_real_yjp36    ;
real dut_real_yjp37    ;
real dut_real_yjp38    ;
real dut_real_yjp39    ;
real dut_real_yjp40    ;
real dut_real_yjp41    ;
real dut_real_yjp42    ;
real dut_real_yjp43    ;
real dut_real_yjp44    ;
real dut_real_yjp45    ;
real dut_real_yjp46    ;
real dut_real_yjp47    ;
real dut_real_yjp48    ;
real dut_real_yjp49    ;
real dut_real_yjp50    ;
real dut_real_yjp51    ;
real dut_real_yjp52    ;
real dut_real_yjp53    ;
real dut_real_yjp54    ;
real dut_real_yjp55    ;
real dut_real_yjp56    ;
real dut_real_yjp57    ;
real dut_real_yjp58    ;
real dut_real_yjp59    ;
real dut_real_yjp60    ;
real dut_real_yjp61    ;
real dut_real_yjp62    ;
real dut_real_yjp63    ;
`endif //ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128
real dut_real_yjp64    ;
real dut_real_yjp65    ;
real dut_real_yjp66    ;
real dut_real_yjp67    ;
real dut_real_yjp68    ;
real dut_real_yjp69    ;
real dut_real_yjp70    ;
real dut_real_yjp71    ;
real dut_real_yjp72    ;
real dut_real_yjp73    ;
real dut_real_yjp74    ;
real dut_real_yjp75    ;
real dut_real_yjp76    ;
real dut_real_yjp77    ;
real dut_real_yjp78    ;
real dut_real_yjp79    ;
real dut_real_yjp80    ;
real dut_real_yjp81    ;
real dut_real_yjp82    ;
real dut_real_yjp83    ;
real dut_real_yjp84    ;
real dut_real_yjp85    ;
real dut_real_yjp86    ;
real dut_real_yjp87    ;
real dut_real_yjp88    ;
real dut_real_yjp89    ;
real dut_real_yjp90    ;
real dut_real_yjp91    ;
real dut_real_yjp92    ;
real dut_real_yjp93    ;
real dut_real_yjp94    ;
real dut_real_yjp95    ;
real dut_real_yjp96    ;
real dut_real_yjp97    ;
real dut_real_yjp98    ;
real dut_real_yjp99    ;
real dut_real_yjp100   ;
real dut_real_yjp101   ;
real dut_real_yjp102   ;
real dut_real_yjp103   ;
real dut_real_yjp104   ;
real dut_real_yjp105   ;
real dut_real_yjp106   ;
real dut_real_yjp107   ;
real dut_real_yjp108   ;
real dut_real_yjp109   ;
real dut_real_yjp110   ;
real dut_real_yjp111   ;
real dut_real_yjp112   ;
real dut_real_yjp113   ;
real dut_real_yjp114   ;
real dut_real_yjp115   ;
real dut_real_yjp116   ;
real dut_real_yjp117   ;
real dut_real_yjp118   ;
real dut_real_yjp119   ;
real dut_real_yjp120   ;
real dut_real_yjp121   ;
real dut_real_yjp122   ;
real dut_real_yjp123   ;
real dut_real_yjp124   ;
real dut_real_yjp125   ;
real dut_real_yjp126   ;
real dut_real_yjp127   ;
`endif //ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256
real dut_real_yjp128   ;
real dut_real_yjp129   ;
real dut_real_yjp130   ;
real dut_real_yjp131   ;
real dut_real_yjp132   ;
real dut_real_yjp133   ;
real dut_real_yjp134   ;
real dut_real_yjp135   ;
real dut_real_yjp136   ;
real dut_real_yjp137   ;
real dut_real_yjp138   ;
real dut_real_yjp139   ;
real dut_real_yjp140   ;
real dut_real_yjp141   ;
real dut_real_yjp142   ;
real dut_real_yjp143   ;
real dut_real_yjp144   ;
real dut_real_yjp145   ;
real dut_real_yjp146   ;
real dut_real_yjp147   ;
real dut_real_yjp148   ;
real dut_real_yjp149   ;
real dut_real_yjp150   ;
real dut_real_yjp151   ;
real dut_real_yjp152   ;
real dut_real_yjp153   ;
real dut_real_yjp154   ;
real dut_real_yjp155   ;
real dut_real_yjp156   ;
real dut_real_yjp157   ;
real dut_real_yjp158   ;
real dut_real_yjp159   ;
real dut_real_yjp160   ;
real dut_real_yjp161   ;
real dut_real_yjp162   ;
real dut_real_yjp163   ;
real dut_real_yjp164   ;
real dut_real_yjp165   ;
real dut_real_yjp166   ;
real dut_real_yjp167   ;
real dut_real_yjp168   ;
real dut_real_yjp169   ;
real dut_real_yjp170   ;
real dut_real_yjp171   ;
real dut_real_yjp172   ;
real dut_real_yjp173   ;
real dut_real_yjp174   ;
real dut_real_yjp175   ;
real dut_real_yjp176   ;
real dut_real_yjp177   ;
real dut_real_yjp178   ;
real dut_real_yjp179   ;
real dut_real_yjp180   ;
real dut_real_yjp181   ;
real dut_real_yjp182   ;
real dut_real_yjp183   ;
real dut_real_yjp184   ;
real dut_real_yjp185   ;
real dut_real_yjp186   ;
real dut_real_yjp187   ;
real dut_real_yjp188   ;
real dut_real_yjp189   ;
real dut_real_yjp190   ;
real dut_real_yjp191   ;
real dut_real_yjp192   ;
real dut_real_yjp193   ;
real dut_real_yjp194   ;
real dut_real_yjp195   ;
real dut_real_yjp196   ;
real dut_real_yjp197   ;
real dut_real_yjp198   ;
real dut_real_yjp199   ;
real dut_real_yjp200   ;
real dut_real_yjp201   ;
real dut_real_yjp202   ;
real dut_real_yjp203   ;
real dut_real_yjp204   ;
real dut_real_yjp205   ;
real dut_real_yjp206   ;
real dut_real_yjp207   ;
real dut_real_yjp208   ;
real dut_real_yjp209   ;
real dut_real_yjp210   ;
real dut_real_yjp211   ;
real dut_real_yjp212   ;
real dut_real_yjp213   ;
real dut_real_yjp214   ;
real dut_real_yjp215   ;
real dut_real_yjp216   ;
real dut_real_yjp217   ;
real dut_real_yjp218   ;
real dut_real_yjp219   ;
real dut_real_yjp220   ;
real dut_real_yjp221   ;
real dut_real_yjp222   ;
real dut_real_yjp223   ;
real dut_real_yjp224   ;
real dut_real_yjp225   ;
real dut_real_yjp226   ;
real dut_real_yjp227   ;
real dut_real_yjp228   ;
real dut_real_yjp229   ;
real dut_real_yjp230   ;
real dut_real_yjp231   ;
real dut_real_yjp232   ;
real dut_real_yjp233   ;
real dut_real_yjp234   ;
real dut_real_yjp235   ;
real dut_real_yjp236   ;
real dut_real_yjp237   ;
real dut_real_yjp238   ;
real dut_real_yjp239   ;
real dut_real_yjp240   ;
real dut_real_yjp241   ;
real dut_real_yjp242   ;
real dut_real_yjp243   ;
real dut_real_yjp244   ;
real dut_real_yjp245   ;
real dut_real_yjp246   ;
real dut_real_yjp247   ;
real dut_real_yjp248   ;
real dut_real_yjp249   ;
real dut_real_yjp250   ;
real dut_real_yjp251   ;
real dut_real_yjp252   ;
real dut_real_yjp253   ;
real dut_real_yjp254   ;
real dut_real_yjp255   ;
`endif //ST_WIDTH_INF_256
`ifdef ST_WIDTH_INF_16
real error_percent0   ;    
real error_percent1   ;    
real error_percent2   ;    
real error_percent3   ;    
real error_percent4   ;    
real error_percent5   ;    
real error_percent6   ;    
real error_percent7   ;    
real error_percent8   ;    
real error_percent9   ;    
real error_percent10  ;    
real error_percent11  ;    
real error_percent12  ;    
real error_percent13  ;    
real error_percent14  ;    
real error_percent15  ;    
`endif //ST_WIDTH_INF_16
`ifdef ST_WIDTH_INF_32
real error_percent16  ;    
real error_percent17  ;    
real error_percent18  ;    
real error_percent19  ;    
real error_percent20  ;    
real error_percent21  ;    
real error_percent22  ;    
real error_percent23  ;    
real error_percent24  ;    
real error_percent25  ;    
real error_percent26  ;    
real error_percent27  ;    
real error_percent28  ;    
real error_percent29  ;    
real error_percent30  ;    
real error_percent31  ;    
`endif //ST_WIDTH_INF_32
`ifdef ST_WIDTH_INF_64
real error_percent32  ;    
real error_percent33  ;    
real error_percent34  ;    
real error_percent35  ;    
real error_percent36  ;    
real error_percent37  ;    
real error_percent38  ;    
real error_percent39  ;    
real error_percent40  ;    
real error_percent41  ;    
real error_percent42  ;    
real error_percent43  ;    
real error_percent44  ;    
real error_percent45  ;    
real error_percent46  ;    
real error_percent47  ;    
real error_percent48  ;    
real error_percent49  ;    
real error_percent50  ;    
real error_percent51  ;    
real error_percent52  ;    
real error_percent53  ;    
real error_percent54  ;    
real error_percent55  ;    
real error_percent56  ;    
real error_percent57  ;    
real error_percent58  ;    
real error_percent59  ;    
real error_percent60  ;    
real error_percent61  ;    
real error_percent62  ;    
real error_percent63  ;    
`endif //ST_WIDTH_INF_64
`ifdef ST_WIDTH_INF_128
real error_percent64  ;    
real error_percent65  ;    
real error_percent66  ;    
real error_percent67  ;    
real error_percent68  ;    
real error_percent69  ;    
real error_percent70  ;    
real error_percent71  ;    
real error_percent72  ;    
real error_percent73  ;    
real error_percent74  ;    
real error_percent75  ;    
real error_percent76  ;    
real error_percent77  ;    
real error_percent78  ;    
real error_percent79  ;    
real error_percent80  ;    
real error_percent81  ;    
real error_percent82  ;    
real error_percent83  ;    
real error_percent84  ;    
real error_percent85  ;    
real error_percent86  ;    
real error_percent87  ;    
real error_percent88  ;    
real error_percent89  ;    
real error_percent90  ;    
real error_percent91  ;    
real error_percent92  ;    
real error_percent93  ;    
real error_percent94  ;    
real error_percent95  ;    
real error_percent96  ;    
real error_percent97  ;    
real error_percent98  ;    
real error_percent99  ;    
real error_percent100 ;    
real error_percent101 ;    
real error_percent102 ;    
real error_percent103 ;    
real error_percent104 ;    
real error_percent105 ;    
real error_percent106 ;    
real error_percent107 ;    
real error_percent108 ;    
real error_percent109 ;    
real error_percent110 ;    
real error_percent111 ;    
real error_percent112 ;    
real error_percent113 ;    
real error_percent114 ;    
real error_percent115 ;    
real error_percent116 ;    
real error_percent117 ;    
real error_percent118 ;    
real error_percent119 ;    
real error_percent120 ;    
real error_percent121 ;    
real error_percent122 ;    
real error_percent123 ;    
real error_percent124 ;    
real error_percent125 ;    
real error_percent126 ;    
real error_percent127 ;    
`endif //ST_WIDTH_INF_128
`ifdef ST_WIDTH_INF_256
real error_percent128 ;
real error_percent129 ;
real error_percent130 ;
real error_percent131 ;
real error_percent132 ;
real error_percent133 ;
real error_percent134 ;
real error_percent135 ;
real error_percent136 ;
real error_percent137 ;
real error_percent138 ;
real error_percent139 ;
real error_percent140 ;
real error_percent141 ;
real error_percent142 ;
real error_percent143 ;
real error_percent144 ;
real error_percent145 ;
real error_percent146 ;
real error_percent147 ;
real error_percent148 ;
real error_percent149 ;
real error_percent150 ;
real error_percent151 ;
real error_percent152 ;
real error_percent153 ;
real error_percent154 ;
real error_percent155 ;
real error_percent156 ;
real error_percent157 ;
real error_percent158 ;
real error_percent159 ;
real error_percent160 ;
real error_percent161 ;
real error_percent162 ;
real error_percent163 ;
real error_percent164 ;
real error_percent165 ;
real error_percent166 ;
real error_percent167 ;
real error_percent168 ;
real error_percent169 ;
real error_percent170 ;
real error_percent171 ;
real error_percent172 ;
real error_percent173 ;
real error_percent174 ;
real error_percent175 ;
real error_percent176 ;
real error_percent177 ;
real error_percent178 ;
real error_percent179 ;
real error_percent180 ;
real error_percent181 ;
real error_percent182 ;
real error_percent183 ;
real error_percent184 ;
real error_percent185 ;
real error_percent186 ;
real error_percent187 ;
real error_percent188 ;
real error_percent189 ;
real error_percent190 ;
real error_percent191 ;
real error_percent192 ;
real error_percent193 ;
real error_percent194 ;
real error_percent195 ;
real error_percent196 ;
real error_percent197 ;
real error_percent198 ;
real error_percent199 ;
real error_percent200 ;
real error_percent201 ;
real error_percent202 ;
real error_percent203 ;
real error_percent204 ;
real error_percent205 ;
real error_percent206 ;
real error_percent207 ;
real error_percent208 ;
real error_percent209 ;
real error_percent210 ;
real error_percent211 ;
real error_percent212 ;
real error_percent213 ;
real error_percent214 ;
real error_percent215 ;
real error_percent216 ;
real error_percent217 ;
real error_percent218 ;
real error_percent219 ;
real error_percent220 ;
real error_percent221 ;
real error_percent222 ;
real error_percent223 ;
real error_percent224 ;
real error_percent225 ;
real error_percent226 ;
real error_percent227 ;
real error_percent228 ;
real error_percent229 ;
real error_percent230 ;
real error_percent231 ;
real error_percent232 ;
real error_percent233 ;
real error_percent234 ;
real error_percent235 ;
real error_percent236 ;
real error_percent237 ;
real error_percent238 ;
real error_percent239 ;
real error_percent240 ;
real error_percent241 ;
real error_percent242 ;
real error_percent243 ;
real error_percent244 ;
real error_percent245 ;
real error_percent246 ;
real error_percent247 ;
real error_percent248 ;
real error_percent249 ;
real error_percent250 ;
real error_percent251 ;
real error_percent252 ;
real error_percent253 ;
real error_percent254 ;
real error_percent255 ;
`endif // ST_WIDTH_INF_256
